// 
// Standard header to adapt well known macros to our needs.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module Rob_1(
  input         clock,
                reset,
                io_enq_valids_0,
                io_enq_valids_1,
                io_enq_valids_2,
  input  [6:0]  io_enq_uops_0_uopc,
  input         io_enq_uops_0_is_rvc,
                io_enq_uops_0_is_br,
                io_enq_uops_0_is_jalr,
  input  [15:0] io_enq_uops_0_br_mask,
  input  [4:0]  io_enq_uops_0_ftq_idx,
  input         io_enq_uops_0_edge_inst,
  input  [5:0]  io_enq_uops_0_pc_lob,
  input  [6:0]  io_enq_uops_0_rob_idx,
                io_enq_uops_0_pdst,
                io_enq_uops_0_stale_pdst,
  input         io_enq_uops_0_exception,
  input  [63:0] io_enq_uops_0_exc_cause,
  input         io_enq_uops_0_is_fence,
                io_enq_uops_0_is_fencei,
                io_enq_uops_0_uses_ldq,
                io_enq_uops_0_uses_stq,
                io_enq_uops_0_is_sys_pc2epc,
                io_enq_uops_0_is_unique,
                io_enq_uops_0_flush_on_commit,
  input  [5:0]  io_enq_uops_0_ldst,
  input         io_enq_uops_0_ldst_val,
  input  [1:0]  io_enq_uops_0_dst_rtype,
  input         io_enq_uops_0_fp_val,
  input  [6:0]  io_enq_uops_1_uopc,
  input         io_enq_uops_1_is_rvc,
                io_enq_uops_1_is_br,
                io_enq_uops_1_is_jalr,
  input  [15:0] io_enq_uops_1_br_mask,
  input  [4:0]  io_enq_uops_1_ftq_idx,
  input         io_enq_uops_1_edge_inst,
  input  [5:0]  io_enq_uops_1_pc_lob,
  input  [6:0]  io_enq_uops_1_rob_idx,
                io_enq_uops_1_pdst,
                io_enq_uops_1_stale_pdst,
  input         io_enq_uops_1_exception,
  input  [63:0] io_enq_uops_1_exc_cause,
  input         io_enq_uops_1_is_fence,
                io_enq_uops_1_is_fencei,
                io_enq_uops_1_uses_ldq,
                io_enq_uops_1_uses_stq,
                io_enq_uops_1_is_sys_pc2epc,
                io_enq_uops_1_is_unique,
                io_enq_uops_1_flush_on_commit,
  input  [5:0]  io_enq_uops_1_ldst,
  input         io_enq_uops_1_ldst_val,
  input  [1:0]  io_enq_uops_1_dst_rtype,
  input         io_enq_uops_1_fp_val,
  input  [6:0]  io_enq_uops_2_uopc,
  input         io_enq_uops_2_is_rvc,
                io_enq_uops_2_is_br,
                io_enq_uops_2_is_jalr,
  input  [15:0] io_enq_uops_2_br_mask,
  input  [4:0]  io_enq_uops_2_ftq_idx,
  input         io_enq_uops_2_edge_inst,
  input  [5:0]  io_enq_uops_2_pc_lob,
  input  [6:0]  io_enq_uops_2_rob_idx,
                io_enq_uops_2_pdst,
                io_enq_uops_2_stale_pdst,
  input         io_enq_uops_2_exception,
  input  [63:0] io_enq_uops_2_exc_cause,
  input         io_enq_uops_2_is_fence,
                io_enq_uops_2_is_fencei,
                io_enq_uops_2_uses_ldq,
                io_enq_uops_2_uses_stq,
                io_enq_uops_2_is_sys_pc2epc,
                io_enq_uops_2_is_unique,
                io_enq_uops_2_flush_on_commit,
  input  [5:0]  io_enq_uops_2_ldst,
  input         io_enq_uops_2_ldst_val,
  input  [1:0]  io_enq_uops_2_dst_rtype,
  input         io_enq_uops_2_fp_val,
                io_enq_partial_stall,
  input  [39:0] io_xcpt_fetch_pc,
  input  [15:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_rob_idx,
  input         io_brupdate_b2_mispredict,
                io_wb_resps_0_valid,
  input  [6:0]  io_wb_resps_0_bits_uop_rob_idx,
                io_wb_resps_0_bits_uop_pdst,
  input         io_wb_resps_0_bits_predicated,
                io_wb_resps_1_valid,
  input  [6:0]  io_wb_resps_1_bits_uop_rob_idx,
                io_wb_resps_1_bits_uop_pdst,
  input         io_wb_resps_2_valid,
  input  [6:0]  io_wb_resps_2_bits_uop_rob_idx,
                io_wb_resps_2_bits_uop_pdst,
  input         io_wb_resps_3_valid,
  input  [6:0]  io_wb_resps_3_bits_uop_rob_idx,
                io_wb_resps_3_bits_uop_pdst,
  input         io_wb_resps_4_valid,
  input  [6:0]  io_wb_resps_4_bits_uop_rob_idx,
                io_wb_resps_4_bits_uop_pdst,
  input         io_wb_resps_4_bits_predicated,
                io_wb_resps_5_valid,
  input  [6:0]  io_wb_resps_5_bits_uop_rob_idx,
                io_wb_resps_5_bits_uop_pdst,
  input         io_lsu_clr_bsy_0_valid,
  input  [6:0]  io_lsu_clr_bsy_0_bits,
  input         io_lsu_clr_bsy_1_valid,
  input  [6:0]  io_lsu_clr_bsy_1_bits,
  input         io_fflags_0_valid,
  input  [6:0]  io_fflags_0_bits_uop_rob_idx,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_1_valid,
  input  [6:0]  io_fflags_1_bits_uop_rob_idx,
  input  [4:0]  io_fflags_1_bits_flags,
  input         io_lxcpt_valid,
  input  [15:0] io_lxcpt_bits_uop_br_mask,
  input  [6:0]  io_lxcpt_bits_uop_rob_idx,
  input  [4:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  input         io_csr_stall,
  output [6:0]  io_rob_tail_idx,
                io_rob_head_idx,
  output        io_commit_valids_0,
                io_commit_valids_1,
                io_commit_valids_2,
                io_commit_arch_valids_0,
                io_commit_arch_valids_1,
                io_commit_arch_valids_2,
  output [4:0]  io_commit_uops_0_ftq_idx,
  output [6:0]  io_commit_uops_0_pdst,
                io_commit_uops_0_stale_pdst,
  output        io_commit_uops_0_is_fencei,
                io_commit_uops_0_uses_ldq,
                io_commit_uops_0_uses_stq,
  output [5:0]  io_commit_uops_0_ldst,
  output        io_commit_uops_0_ldst_val,
  output [1:0]  io_commit_uops_0_dst_rtype,
  output [4:0]  io_commit_uops_1_ftq_idx,
  output [6:0]  io_commit_uops_1_pdst,
                io_commit_uops_1_stale_pdst,
  output        io_commit_uops_1_is_fencei,
                io_commit_uops_1_uses_ldq,
                io_commit_uops_1_uses_stq,
  output [5:0]  io_commit_uops_1_ldst,
  output        io_commit_uops_1_ldst_val,
  output [1:0]  io_commit_uops_1_dst_rtype,
  output [4:0]  io_commit_uops_2_ftq_idx,
  output [6:0]  io_commit_uops_2_pdst,
                io_commit_uops_2_stale_pdst,
  output        io_commit_uops_2_is_fencei,
                io_commit_uops_2_uses_ldq,
                io_commit_uops_2_uses_stq,
  output [5:0]  io_commit_uops_2_ldst,
  output        io_commit_uops_2_ldst_val,
  output [1:0]  io_commit_uops_2_dst_rtype,
  output        io_commit_fflags_valid,
  output [4:0]  io_commit_fflags_bits,
  output        io_commit_rbk_valids_0,
                io_commit_rbk_valids_1,
                io_commit_rbk_valids_2,
                io_commit_rollback,
                io_com_load_is_at_rob_head,
                io_com_xcpt_valid,
  output [4:0]  io_com_xcpt_bits_ftq_idx,
  output        io_com_xcpt_bits_edge_inst,
  output [5:0]  io_com_xcpt_bits_pc_lob,
  output [63:0] io_com_xcpt_bits_cause,
                io_com_xcpt_bits_badvaddr,
  output        io_flush_valid,
  output [4:0]  io_flush_bits_ftq_idx,
  output        io_flush_bits_edge_inst,
                io_flush_bits_is_rvc,
  output [5:0]  io_flush_bits_pc_lob,
  output [2:0]  io_flush_bits_flush_typ,
  output        io_empty,
                io_ready,
                io_flush_frontend
);

  wire             empty;	// rob.scala:788:41
  wire             full;	// rob.scala:787:39
  wire             will_commit_2;	// rob.scala:547:70
  wire             will_commit_1;	// rob.scala:547:70
  wire             will_commit_0;	// rob.scala:547:70
  wire [4:0]       _rob_fflags_2_ext_R0_data;	// rob.scala:313:28
  wire [4:0]       _rob_fflags_1_ext_R0_data;	// rob.scala:313:28
  wire [4:0]       _rob_fflags_ext_R0_data;	// rob.scala:313:28
  reg  [1:0]       rob_state;	// rob.scala:221:26
  reg  [4:0]       rob_head;	// rob.scala:224:29
  reg  [1:0]       rob_head_lsb;	// rob.scala:225:29
  wire [6:0]       rob_head_idx = {rob_head, rob_head_lsb};	// Cat.scala:30:58, rob.scala:224:29, :225:29
  reg  [4:0]       rob_tail;	// rob.scala:228:29
  reg  [1:0]       rob_tail_lsb;	// rob.scala:229:29
  wire [6:0]       rob_tail_idx = {rob_tail, rob_tail_lsb};	// Cat.scala:30:58, rob.scala:228:29, :229:29
  reg  [4:0]       rob_pnr;	// rob.scala:232:29
  reg  [1:0]       rob_pnr_lsb;	// rob.scala:233:29
  wire             _io_commit_rollback_T_2 = rob_state == 2'h2;	// rob.scala:221:26, :236:31
  wire [4:0]       com_idx = _io_commit_rollback_T_2 ? rob_tail : rob_head;	// rob.scala:224:29, :228:29, :236:{20,31}
  reg              maybe_full;	// rob.scala:239:29
  reg              r_xcpt_val;	// rob.scala:258:33
  reg  [15:0]      r_xcpt_uop_br_mask;	// rob.scala:259:29
  reg  [6:0]       r_xcpt_uop_rob_idx;	// rob.scala:259:29
  reg  [63:0]      r_xcpt_uop_exc_cause;	// rob.scala:259:29
  reg  [39:0]      r_xcpt_badvaddr;	// rob.scala:260:29
  reg              rob_val_0;	// rob.scala:307:32
  reg              rob_val_1;	// rob.scala:307:32
  reg              rob_val_2;	// rob.scala:307:32
  reg              rob_val_3;	// rob.scala:307:32
  reg              rob_val_4;	// rob.scala:307:32
  reg              rob_val_5;	// rob.scala:307:32
  reg              rob_val_6;	// rob.scala:307:32
  reg              rob_val_7;	// rob.scala:307:32
  reg              rob_val_8;	// rob.scala:307:32
  reg              rob_val_9;	// rob.scala:307:32
  reg              rob_val_10;	// rob.scala:307:32
  reg              rob_val_11;	// rob.scala:307:32
  reg              rob_val_12;	// rob.scala:307:32
  reg              rob_val_13;	// rob.scala:307:32
  reg              rob_val_14;	// rob.scala:307:32
  reg              rob_val_15;	// rob.scala:307:32
  reg              rob_val_16;	// rob.scala:307:32
  reg              rob_val_17;	// rob.scala:307:32
  reg              rob_val_18;	// rob.scala:307:32
  reg              rob_val_19;	// rob.scala:307:32
  reg              rob_val_20;	// rob.scala:307:32
  reg              rob_val_21;	// rob.scala:307:32
  reg              rob_val_22;	// rob.scala:307:32
  reg              rob_val_23;	// rob.scala:307:32
  reg              rob_val_24;	// rob.scala:307:32
  reg              rob_val_25;	// rob.scala:307:32
  reg              rob_val_26;	// rob.scala:307:32
  reg              rob_val_27;	// rob.scala:307:32
  reg              rob_val_28;	// rob.scala:307:32
  reg              rob_val_29;	// rob.scala:307:32
  reg              rob_val_30;	// rob.scala:307:32
  reg              rob_val_31;	// rob.scala:307:32
  reg              rob_bsy_0;	// rob.scala:308:28
  reg              rob_bsy_1;	// rob.scala:308:28
  reg              rob_bsy_2;	// rob.scala:308:28
  reg              rob_bsy_3;	// rob.scala:308:28
  reg              rob_bsy_4;	// rob.scala:308:28
  reg              rob_bsy_5;	// rob.scala:308:28
  reg              rob_bsy_6;	// rob.scala:308:28
  reg              rob_bsy_7;	// rob.scala:308:28
  reg              rob_bsy_8;	// rob.scala:308:28
  reg              rob_bsy_9;	// rob.scala:308:28
  reg              rob_bsy_10;	// rob.scala:308:28
  reg              rob_bsy_11;	// rob.scala:308:28
  reg              rob_bsy_12;	// rob.scala:308:28
  reg              rob_bsy_13;	// rob.scala:308:28
  reg              rob_bsy_14;	// rob.scala:308:28
  reg              rob_bsy_15;	// rob.scala:308:28
  reg              rob_bsy_16;	// rob.scala:308:28
  reg              rob_bsy_17;	// rob.scala:308:28
  reg              rob_bsy_18;	// rob.scala:308:28
  reg              rob_bsy_19;	// rob.scala:308:28
  reg              rob_bsy_20;	// rob.scala:308:28
  reg              rob_bsy_21;	// rob.scala:308:28
  reg              rob_bsy_22;	// rob.scala:308:28
  reg              rob_bsy_23;	// rob.scala:308:28
  reg              rob_bsy_24;	// rob.scala:308:28
  reg              rob_bsy_25;	// rob.scala:308:28
  reg              rob_bsy_26;	// rob.scala:308:28
  reg              rob_bsy_27;	// rob.scala:308:28
  reg              rob_bsy_28;	// rob.scala:308:28
  reg              rob_bsy_29;	// rob.scala:308:28
  reg              rob_bsy_30;	// rob.scala:308:28
  reg              rob_bsy_31;	// rob.scala:308:28
  reg              rob_unsafe_0;	// rob.scala:309:28
  reg              rob_unsafe_1;	// rob.scala:309:28
  reg              rob_unsafe_2;	// rob.scala:309:28
  reg              rob_unsafe_3;	// rob.scala:309:28
  reg              rob_unsafe_4;	// rob.scala:309:28
  reg              rob_unsafe_5;	// rob.scala:309:28
  reg              rob_unsafe_6;	// rob.scala:309:28
  reg              rob_unsafe_7;	// rob.scala:309:28
  reg              rob_unsafe_8;	// rob.scala:309:28
  reg              rob_unsafe_9;	// rob.scala:309:28
  reg              rob_unsafe_10;	// rob.scala:309:28
  reg              rob_unsafe_11;	// rob.scala:309:28
  reg              rob_unsafe_12;	// rob.scala:309:28
  reg              rob_unsafe_13;	// rob.scala:309:28
  reg              rob_unsafe_14;	// rob.scala:309:28
  reg              rob_unsafe_15;	// rob.scala:309:28
  reg              rob_unsafe_16;	// rob.scala:309:28
  reg              rob_unsafe_17;	// rob.scala:309:28
  reg              rob_unsafe_18;	// rob.scala:309:28
  reg              rob_unsafe_19;	// rob.scala:309:28
  reg              rob_unsafe_20;	// rob.scala:309:28
  reg              rob_unsafe_21;	// rob.scala:309:28
  reg              rob_unsafe_22;	// rob.scala:309:28
  reg              rob_unsafe_23;	// rob.scala:309:28
  reg              rob_unsafe_24;	// rob.scala:309:28
  reg              rob_unsafe_25;	// rob.scala:309:28
  reg              rob_unsafe_26;	// rob.scala:309:28
  reg              rob_unsafe_27;	// rob.scala:309:28
  reg              rob_unsafe_28;	// rob.scala:309:28
  reg              rob_unsafe_29;	// rob.scala:309:28
  reg              rob_unsafe_30;	// rob.scala:309:28
  reg              rob_unsafe_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_0_uopc;	// rob.scala:310:28
  reg              rob_uop_0_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_0_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_0_ldst;	// rob.scala:310:28
  reg              rob_uop_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_uopc;	// rob.scala:310:28
  reg              rob_uop_1_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_ldst;	// rob.scala:310:28
  reg              rob_uop_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_uopc;	// rob.scala:310:28
  reg              rob_uop_2_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_ldst;	// rob.scala:310:28
  reg              rob_uop_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_uopc;	// rob.scala:310:28
  reg              rob_uop_3_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_3_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_3_ldst;	// rob.scala:310:28
  reg              rob_uop_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_4_uopc;	// rob.scala:310:28
  reg              rob_uop_4_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_4_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_4_ldst;	// rob.scala:310:28
  reg              rob_uop_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_5_uopc;	// rob.scala:310:28
  reg              rob_uop_5_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_5_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_5_ldst;	// rob.scala:310:28
  reg              rob_uop_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_6_uopc;	// rob.scala:310:28
  reg              rob_uop_6_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_6_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_6_ldst;	// rob.scala:310:28
  reg              rob_uop_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_7_uopc;	// rob.scala:310:28
  reg              rob_uop_7_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_7_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_7_ldst;	// rob.scala:310:28
  reg              rob_uop_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_8_uopc;	// rob.scala:310:28
  reg              rob_uop_8_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_8_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_8_ldst;	// rob.scala:310:28
  reg              rob_uop_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_9_uopc;	// rob.scala:310:28
  reg              rob_uop_9_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_9_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_9_ldst;	// rob.scala:310:28
  reg              rob_uop_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_10_uopc;	// rob.scala:310:28
  reg              rob_uop_10_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_10_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_10_ldst;	// rob.scala:310:28
  reg              rob_uop_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_11_uopc;	// rob.scala:310:28
  reg              rob_uop_11_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_11_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_11_ldst;	// rob.scala:310:28
  reg              rob_uop_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_12_uopc;	// rob.scala:310:28
  reg              rob_uop_12_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_12_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_12_ldst;	// rob.scala:310:28
  reg              rob_uop_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_13_uopc;	// rob.scala:310:28
  reg              rob_uop_13_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_13_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_13_ldst;	// rob.scala:310:28
  reg              rob_uop_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_14_uopc;	// rob.scala:310:28
  reg              rob_uop_14_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_14_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_14_ldst;	// rob.scala:310:28
  reg              rob_uop_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_15_uopc;	// rob.scala:310:28
  reg              rob_uop_15_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_15_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_15_ldst;	// rob.scala:310:28
  reg              rob_uop_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_16_uopc;	// rob.scala:310:28
  reg              rob_uop_16_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_16_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_16_ldst;	// rob.scala:310:28
  reg              rob_uop_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_17_uopc;	// rob.scala:310:28
  reg              rob_uop_17_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_17_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_17_ldst;	// rob.scala:310:28
  reg              rob_uop_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_18_uopc;	// rob.scala:310:28
  reg              rob_uop_18_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_18_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_18_ldst;	// rob.scala:310:28
  reg              rob_uop_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_19_uopc;	// rob.scala:310:28
  reg              rob_uop_19_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_19_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_19_ldst;	// rob.scala:310:28
  reg              rob_uop_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_20_uopc;	// rob.scala:310:28
  reg              rob_uop_20_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_20_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_20_ldst;	// rob.scala:310:28
  reg              rob_uop_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_21_uopc;	// rob.scala:310:28
  reg              rob_uop_21_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_21_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_21_ldst;	// rob.scala:310:28
  reg              rob_uop_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_22_uopc;	// rob.scala:310:28
  reg              rob_uop_22_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_22_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_22_ldst;	// rob.scala:310:28
  reg              rob_uop_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_23_uopc;	// rob.scala:310:28
  reg              rob_uop_23_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_23_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_23_ldst;	// rob.scala:310:28
  reg              rob_uop_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_24_uopc;	// rob.scala:310:28
  reg              rob_uop_24_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_24_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_24_ldst;	// rob.scala:310:28
  reg              rob_uop_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_25_uopc;	// rob.scala:310:28
  reg              rob_uop_25_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_25_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_25_ldst;	// rob.scala:310:28
  reg              rob_uop_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_26_uopc;	// rob.scala:310:28
  reg              rob_uop_26_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_26_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_26_ldst;	// rob.scala:310:28
  reg              rob_uop_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_27_uopc;	// rob.scala:310:28
  reg              rob_uop_27_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_27_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_27_ldst;	// rob.scala:310:28
  reg              rob_uop_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_28_uopc;	// rob.scala:310:28
  reg              rob_uop_28_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_28_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_28_ldst;	// rob.scala:310:28
  reg              rob_uop_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_29_uopc;	// rob.scala:310:28
  reg              rob_uop_29_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_29_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_29_ldst;	// rob.scala:310:28
  reg              rob_uop_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_30_uopc;	// rob.scala:310:28
  reg              rob_uop_30_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_30_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_30_ldst;	// rob.scala:310:28
  reg              rob_uop_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_31_uopc;	// rob.scala:310:28
  reg              rob_uop_31_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_31_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_31_ldst;	// rob.scala:310:28
  reg              rob_uop_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_0;	// rob.scala:311:28
  reg              rob_exception_1;	// rob.scala:311:28
  reg              rob_exception_2;	// rob.scala:311:28
  reg              rob_exception_3;	// rob.scala:311:28
  reg              rob_exception_4;	// rob.scala:311:28
  reg              rob_exception_5;	// rob.scala:311:28
  reg              rob_exception_6;	// rob.scala:311:28
  reg              rob_exception_7;	// rob.scala:311:28
  reg              rob_exception_8;	// rob.scala:311:28
  reg              rob_exception_9;	// rob.scala:311:28
  reg              rob_exception_10;	// rob.scala:311:28
  reg              rob_exception_11;	// rob.scala:311:28
  reg              rob_exception_12;	// rob.scala:311:28
  reg              rob_exception_13;	// rob.scala:311:28
  reg              rob_exception_14;	// rob.scala:311:28
  reg              rob_exception_15;	// rob.scala:311:28
  reg              rob_exception_16;	// rob.scala:311:28
  reg              rob_exception_17;	// rob.scala:311:28
  reg              rob_exception_18;	// rob.scala:311:28
  reg              rob_exception_19;	// rob.scala:311:28
  reg              rob_exception_20;	// rob.scala:311:28
  reg              rob_exception_21;	// rob.scala:311:28
  reg              rob_exception_22;	// rob.scala:311:28
  reg              rob_exception_23;	// rob.scala:311:28
  reg              rob_exception_24;	// rob.scala:311:28
  reg              rob_exception_25;	// rob.scala:311:28
  reg              rob_exception_26;	// rob.scala:311:28
  reg              rob_exception_27;	// rob.scala:311:28
  reg              rob_exception_28;	// rob.scala:311:28
  reg              rob_exception_29;	// rob.scala:311:28
  reg              rob_exception_30;	// rob.scala:311:28
  reg              rob_exception_31;	// rob.scala:311:28
  reg              rob_predicated_0;	// rob.scala:312:29
  reg              rob_predicated_1;	// rob.scala:312:29
  reg              rob_predicated_2;	// rob.scala:312:29
  reg              rob_predicated_3;	// rob.scala:312:29
  reg              rob_predicated_4;	// rob.scala:312:29
  reg              rob_predicated_5;	// rob.scala:312:29
  reg              rob_predicated_6;	// rob.scala:312:29
  reg              rob_predicated_7;	// rob.scala:312:29
  reg              rob_predicated_8;	// rob.scala:312:29
  reg              rob_predicated_9;	// rob.scala:312:29
  reg              rob_predicated_10;	// rob.scala:312:29
  reg              rob_predicated_11;	// rob.scala:312:29
  reg              rob_predicated_12;	// rob.scala:312:29
  reg              rob_predicated_13;	// rob.scala:312:29
  reg              rob_predicated_14;	// rob.scala:312:29
  reg              rob_predicated_15;	// rob.scala:312:29
  reg              rob_predicated_16;	// rob.scala:312:29
  reg              rob_predicated_17;	// rob.scala:312:29
  reg              rob_predicated_18;	// rob.scala:312:29
  reg              rob_predicated_19;	// rob.scala:312:29
  reg              rob_predicated_20;	// rob.scala:312:29
  reg              rob_predicated_21;	// rob.scala:312:29
  reg              rob_predicated_22;	// rob.scala:312:29
  reg              rob_predicated_23;	// rob.scala:312:29
  reg              rob_predicated_24;	// rob.scala:312:29
  reg              rob_predicated_25;	// rob.scala:312:29
  reg              rob_predicated_26;	// rob.scala:312:29
  reg              rob_predicated_27;	// rob.scala:312:29
  reg              rob_predicated_28;	// rob.scala:312:29
  reg              rob_predicated_29;	// rob.scala:312:29
  reg              rob_predicated_30;	// rob.scala:312:29
  reg              rob_predicated_31;	// rob.scala:312:29
  wire [31:0]      _GEN =
    {{rob_val_31},
     {rob_val_30},
     {rob_val_29},
     {rob_val_28},
     {rob_val_27},
     {rob_val_26},
     {rob_val_25},
     {rob_val_24},
     {rob_val_23},
     {rob_val_22},
     {rob_val_21},
     {rob_val_20},
     {rob_val_19},
     {rob_val_18},
     {rob_val_17},
     {rob_val_16},
     {rob_val_15},
     {rob_val_14},
     {rob_val_13},
     {rob_val_12},
     {rob_val_11},
     {rob_val_10},
     {rob_val_9},
     {rob_val_8},
     {rob_val_7},
     {rob_val_6},
     {rob_val_5},
     {rob_val_4},
     {rob_val_3},
     {rob_val_2},
     {rob_val_1},
     {rob_val_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_0 = _GEN[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_0 =
    io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_1 =
    io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_2 =
    io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_3 =
    io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_4 =
    io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_5 =
    io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :346:27
  wire             _GEN_6 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :361:31
  wire [31:0]      _GEN_7 =
    {{rob_bsy_31},
     {rob_bsy_30},
     {rob_bsy_29},
     {rob_bsy_28},
     {rob_bsy_27},
     {rob_bsy_26},
     {rob_bsy_25},
     {rob_bsy_24},
     {rob_bsy_23},
     {rob_bsy_22},
     {rob_bsy_21},
     {rob_bsy_20},
     {rob_bsy_19},
     {rob_bsy_18},
     {rob_bsy_17},
     {rob_bsy_16},
     {rob_bsy_15},
     {rob_bsy_14},
     {rob_bsy_13},
     {rob_bsy_12},
     {rob_bsy_11},
     {rob_bsy_10},
     {rob_bsy_9},
     {rob_bsy_8},
     {rob_bsy_7},
     {rob_bsy_6},
     {rob_bsy_5},
     {rob_bsy_4},
     {rob_bsy_3},
     {rob_bsy_2},
     {rob_bsy_1},
     {rob_bsy_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_8 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :361:31
  wire             _GEN_9 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h0;	// rob.scala:221:26, :272:36, :304:53, :390:26
  wire [31:0]      _GEN_10 =
    {{rob_unsafe_31},
     {rob_unsafe_30},
     {rob_unsafe_29},
     {rob_unsafe_28},
     {rob_unsafe_27},
     {rob_unsafe_26},
     {rob_unsafe_25},
     {rob_unsafe_24},
     {rob_unsafe_23},
     {rob_unsafe_22},
     {rob_unsafe_21},
     {rob_unsafe_20},
     {rob_unsafe_19},
     {rob_unsafe_18},
     {rob_unsafe_17},
     {rob_unsafe_16},
     {rob_unsafe_15},
     {rob_unsafe_14},
     {rob_unsafe_13},
     {rob_unsafe_12},
     {rob_unsafe_11},
     {rob_unsafe_10},
     {rob_unsafe_9},
     {rob_unsafe_8},
     {rob_unsafe_7},
     {rob_unsafe_6},
     {rob_unsafe_5},
     {rob_unsafe_4},
     {rob_unsafe_3},
     {rob_unsafe_2},
     {rob_unsafe_1},
     {rob_unsafe_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_0 = _GEN[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_11 =
    {{rob_exception_31},
     {rob_exception_30},
     {rob_exception_29},
     {rob_exception_28},
     {rob_exception_27},
     {rob_exception_26},
     {rob_exception_25},
     {rob_exception_24},
     {rob_exception_23},
     {rob_exception_22},
     {rob_exception_21},
     {rob_exception_20},
     {rob_exception_19},
     {rob_exception_18},
     {rob_exception_17},
     {rob_exception_16},
     {rob_exception_15},
     {rob_exception_14},
     {rob_exception_13},
     {rob_exception_12},
     {rob_exception_11},
     {rob_exception_10},
     {rob_exception_9},
     {rob_exception_8},
     {rob_exception_7},
     {rob_exception_6},
     {rob_exception_5},
     {rob_exception_4},
     {rob_exception_3},
     {rob_exception_2},
     {rob_exception_1},
     {rob_exception_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_0 = rob_head_vals_0 & _GEN_11[rob_head];	// rob.scala:224:29, :398:49
  wire             can_commit_0 = rob_head_vals_0 & ~_GEN_7[rob_head] & ~io_csr_stall;	// rob.scala:224:29, :366:31, :398:49, :404:{43,64,67}
  wire [31:0]      _GEN_12 =
    {{rob_predicated_31},
     {rob_predicated_30},
     {rob_predicated_29},
     {rob_predicated_28},
     {rob_predicated_27},
     {rob_predicated_26},
     {rob_predicated_25},
     {rob_predicated_24},
     {rob_predicated_23},
     {rob_predicated_22},
     {rob_predicated_21},
     {rob_predicated_20},
     {rob_predicated_19},
     {rob_predicated_18},
     {rob_predicated_17},
     {rob_predicated_16},
     {rob_predicated_15},
     {rob_predicated_14},
     {rob_predicated_13},
     {rob_predicated_12},
     {rob_predicated_11},
     {rob_predicated_10},
     {rob_predicated_9},
     {rob_predicated_8},
     {rob_predicated_7},
     {rob_predicated_6},
     {rob_predicated_5},
     {rob_predicated_4},
     {rob_predicated_3},
     {rob_predicated_2},
     {rob_predicated_1},
     {rob_predicated_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_13 =
    {{rob_uop_31_uopc},
     {rob_uop_30_uopc},
     {rob_uop_29_uopc},
     {rob_uop_28_uopc},
     {rob_uop_27_uopc},
     {rob_uop_26_uopc},
     {rob_uop_25_uopc},
     {rob_uop_24_uopc},
     {rob_uop_23_uopc},
     {rob_uop_22_uopc},
     {rob_uop_21_uopc},
     {rob_uop_20_uopc},
     {rob_uop_19_uopc},
     {rob_uop_18_uopc},
     {rob_uop_17_uopc},
     {rob_uop_16_uopc},
     {rob_uop_15_uopc},
     {rob_uop_14_uopc},
     {rob_uop_13_uopc},
     {rob_uop_12_uopc},
     {rob_uop_11_uopc},
     {rob_uop_10_uopc},
     {rob_uop_9_uopc},
     {rob_uop_8_uopc},
     {rob_uop_7_uopc},
     {rob_uop_6_uopc},
     {rob_uop_5_uopc},
     {rob_uop_4_uopc},
     {rob_uop_3_uopc},
     {rob_uop_2_uopc},
     {rob_uop_1_uopc},
     {rob_uop_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_14 =
    {{rob_uop_31_is_rvc},
     {rob_uop_30_is_rvc},
     {rob_uop_29_is_rvc},
     {rob_uop_28_is_rvc},
     {rob_uop_27_is_rvc},
     {rob_uop_26_is_rvc},
     {rob_uop_25_is_rvc},
     {rob_uop_24_is_rvc},
     {rob_uop_23_is_rvc},
     {rob_uop_22_is_rvc},
     {rob_uop_21_is_rvc},
     {rob_uop_20_is_rvc},
     {rob_uop_19_is_rvc},
     {rob_uop_18_is_rvc},
     {rob_uop_17_is_rvc},
     {rob_uop_16_is_rvc},
     {rob_uop_15_is_rvc},
     {rob_uop_14_is_rvc},
     {rob_uop_13_is_rvc},
     {rob_uop_12_is_rvc},
     {rob_uop_11_is_rvc},
     {rob_uop_10_is_rvc},
     {rob_uop_9_is_rvc},
     {rob_uop_8_is_rvc},
     {rob_uop_7_is_rvc},
     {rob_uop_6_is_rvc},
     {rob_uop_5_is_rvc},
     {rob_uop_4_is_rvc},
     {rob_uop_3_is_rvc},
     {rob_uop_2_is_rvc},
     {rob_uop_1_is_rvc},
     {rob_uop_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][4:0] _GEN_15 =
    {{rob_uop_31_ftq_idx},
     {rob_uop_30_ftq_idx},
     {rob_uop_29_ftq_idx},
     {rob_uop_28_ftq_idx},
     {rob_uop_27_ftq_idx},
     {rob_uop_26_ftq_idx},
     {rob_uop_25_ftq_idx},
     {rob_uop_24_ftq_idx},
     {rob_uop_23_ftq_idx},
     {rob_uop_22_ftq_idx},
     {rob_uop_21_ftq_idx},
     {rob_uop_20_ftq_idx},
     {rob_uop_19_ftq_idx},
     {rob_uop_18_ftq_idx},
     {rob_uop_17_ftq_idx},
     {rob_uop_16_ftq_idx},
     {rob_uop_15_ftq_idx},
     {rob_uop_14_ftq_idx},
     {rob_uop_13_ftq_idx},
     {rob_uop_12_ftq_idx},
     {rob_uop_11_ftq_idx},
     {rob_uop_10_ftq_idx},
     {rob_uop_9_ftq_idx},
     {rob_uop_8_ftq_idx},
     {rob_uop_7_ftq_idx},
     {rob_uop_6_ftq_idx},
     {rob_uop_5_ftq_idx},
     {rob_uop_4_ftq_idx},
     {rob_uop_3_ftq_idx},
     {rob_uop_2_ftq_idx},
     {rob_uop_1_ftq_idx},
     {rob_uop_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_16 =
    {{rob_uop_31_edge_inst},
     {rob_uop_30_edge_inst},
     {rob_uop_29_edge_inst},
     {rob_uop_28_edge_inst},
     {rob_uop_27_edge_inst},
     {rob_uop_26_edge_inst},
     {rob_uop_25_edge_inst},
     {rob_uop_24_edge_inst},
     {rob_uop_23_edge_inst},
     {rob_uop_22_edge_inst},
     {rob_uop_21_edge_inst},
     {rob_uop_20_edge_inst},
     {rob_uop_19_edge_inst},
     {rob_uop_18_edge_inst},
     {rob_uop_17_edge_inst},
     {rob_uop_16_edge_inst},
     {rob_uop_15_edge_inst},
     {rob_uop_14_edge_inst},
     {rob_uop_13_edge_inst},
     {rob_uop_12_edge_inst},
     {rob_uop_11_edge_inst},
     {rob_uop_10_edge_inst},
     {rob_uop_9_edge_inst},
     {rob_uop_8_edge_inst},
     {rob_uop_7_edge_inst},
     {rob_uop_6_edge_inst},
     {rob_uop_5_edge_inst},
     {rob_uop_4_edge_inst},
     {rob_uop_3_edge_inst},
     {rob_uop_2_edge_inst},
     {rob_uop_1_edge_inst},
     {rob_uop_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_17 =
    {{rob_uop_31_pc_lob},
     {rob_uop_30_pc_lob},
     {rob_uop_29_pc_lob},
     {rob_uop_28_pc_lob},
     {rob_uop_27_pc_lob},
     {rob_uop_26_pc_lob},
     {rob_uop_25_pc_lob},
     {rob_uop_24_pc_lob},
     {rob_uop_23_pc_lob},
     {rob_uop_22_pc_lob},
     {rob_uop_21_pc_lob},
     {rob_uop_20_pc_lob},
     {rob_uop_19_pc_lob},
     {rob_uop_18_pc_lob},
     {rob_uop_17_pc_lob},
     {rob_uop_16_pc_lob},
     {rob_uop_15_pc_lob},
     {rob_uop_14_pc_lob},
     {rob_uop_13_pc_lob},
     {rob_uop_12_pc_lob},
     {rob_uop_11_pc_lob},
     {rob_uop_10_pc_lob},
     {rob_uop_9_pc_lob},
     {rob_uop_8_pc_lob},
     {rob_uop_7_pc_lob},
     {rob_uop_6_pc_lob},
     {rob_uop_5_pc_lob},
     {rob_uop_4_pc_lob},
     {rob_uop_3_pc_lob},
     {rob_uop_2_pc_lob},
     {rob_uop_1_pc_lob},
     {rob_uop_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_18 =
    {{rob_uop_31_pdst},
     {rob_uop_30_pdst},
     {rob_uop_29_pdst},
     {rob_uop_28_pdst},
     {rob_uop_27_pdst},
     {rob_uop_26_pdst},
     {rob_uop_25_pdst},
     {rob_uop_24_pdst},
     {rob_uop_23_pdst},
     {rob_uop_22_pdst},
     {rob_uop_21_pdst},
     {rob_uop_20_pdst},
     {rob_uop_19_pdst},
     {rob_uop_18_pdst},
     {rob_uop_17_pdst},
     {rob_uop_16_pdst},
     {rob_uop_15_pdst},
     {rob_uop_14_pdst},
     {rob_uop_13_pdst},
     {rob_uop_12_pdst},
     {rob_uop_11_pdst},
     {rob_uop_10_pdst},
     {rob_uop_9_pdst},
     {rob_uop_8_pdst},
     {rob_uop_7_pdst},
     {rob_uop_6_pdst},
     {rob_uop_5_pdst},
     {rob_uop_4_pdst},
     {rob_uop_3_pdst},
     {rob_uop_2_pdst},
     {rob_uop_1_pdst},
     {rob_uop_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_19 =
    {{rob_uop_31_stale_pdst},
     {rob_uop_30_stale_pdst},
     {rob_uop_29_stale_pdst},
     {rob_uop_28_stale_pdst},
     {rob_uop_27_stale_pdst},
     {rob_uop_26_stale_pdst},
     {rob_uop_25_stale_pdst},
     {rob_uop_24_stale_pdst},
     {rob_uop_23_stale_pdst},
     {rob_uop_22_stale_pdst},
     {rob_uop_21_stale_pdst},
     {rob_uop_20_stale_pdst},
     {rob_uop_19_stale_pdst},
     {rob_uop_18_stale_pdst},
     {rob_uop_17_stale_pdst},
     {rob_uop_16_stale_pdst},
     {rob_uop_15_stale_pdst},
     {rob_uop_14_stale_pdst},
     {rob_uop_13_stale_pdst},
     {rob_uop_12_stale_pdst},
     {rob_uop_11_stale_pdst},
     {rob_uop_10_stale_pdst},
     {rob_uop_9_stale_pdst},
     {rob_uop_8_stale_pdst},
     {rob_uop_7_stale_pdst},
     {rob_uop_6_stale_pdst},
     {rob_uop_5_stale_pdst},
     {rob_uop_4_stale_pdst},
     {rob_uop_3_stale_pdst},
     {rob_uop_2_stale_pdst},
     {rob_uop_1_stale_pdst},
     {rob_uop_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_20 =
    {{rob_uop_31_is_fencei},
     {rob_uop_30_is_fencei},
     {rob_uop_29_is_fencei},
     {rob_uop_28_is_fencei},
     {rob_uop_27_is_fencei},
     {rob_uop_26_is_fencei},
     {rob_uop_25_is_fencei},
     {rob_uop_24_is_fencei},
     {rob_uop_23_is_fencei},
     {rob_uop_22_is_fencei},
     {rob_uop_21_is_fencei},
     {rob_uop_20_is_fencei},
     {rob_uop_19_is_fencei},
     {rob_uop_18_is_fencei},
     {rob_uop_17_is_fencei},
     {rob_uop_16_is_fencei},
     {rob_uop_15_is_fencei},
     {rob_uop_14_is_fencei},
     {rob_uop_13_is_fencei},
     {rob_uop_12_is_fencei},
     {rob_uop_11_is_fencei},
     {rob_uop_10_is_fencei},
     {rob_uop_9_is_fencei},
     {rob_uop_8_is_fencei},
     {rob_uop_7_is_fencei},
     {rob_uop_6_is_fencei},
     {rob_uop_5_is_fencei},
     {rob_uop_4_is_fencei},
     {rob_uop_3_is_fencei},
     {rob_uop_2_is_fencei},
     {rob_uop_1_is_fencei},
     {rob_uop_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_21 =
    {{rob_uop_31_uses_ldq},
     {rob_uop_30_uses_ldq},
     {rob_uop_29_uses_ldq},
     {rob_uop_28_uses_ldq},
     {rob_uop_27_uses_ldq},
     {rob_uop_26_uses_ldq},
     {rob_uop_25_uses_ldq},
     {rob_uop_24_uses_ldq},
     {rob_uop_23_uses_ldq},
     {rob_uop_22_uses_ldq},
     {rob_uop_21_uses_ldq},
     {rob_uop_20_uses_ldq},
     {rob_uop_19_uses_ldq},
     {rob_uop_18_uses_ldq},
     {rob_uop_17_uses_ldq},
     {rob_uop_16_uses_ldq},
     {rob_uop_15_uses_ldq},
     {rob_uop_14_uses_ldq},
     {rob_uop_13_uses_ldq},
     {rob_uop_12_uses_ldq},
     {rob_uop_11_uses_ldq},
     {rob_uop_10_uses_ldq},
     {rob_uop_9_uses_ldq},
     {rob_uop_8_uses_ldq},
     {rob_uop_7_uses_ldq},
     {rob_uop_6_uses_ldq},
     {rob_uop_5_uses_ldq},
     {rob_uop_4_uses_ldq},
     {rob_uop_3_uses_ldq},
     {rob_uop_2_uses_ldq},
     {rob_uop_1_uses_ldq},
     {rob_uop_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_22 =
    {{rob_uop_31_uses_stq},
     {rob_uop_30_uses_stq},
     {rob_uop_29_uses_stq},
     {rob_uop_28_uses_stq},
     {rob_uop_27_uses_stq},
     {rob_uop_26_uses_stq},
     {rob_uop_25_uses_stq},
     {rob_uop_24_uses_stq},
     {rob_uop_23_uses_stq},
     {rob_uop_22_uses_stq},
     {rob_uop_21_uses_stq},
     {rob_uop_20_uses_stq},
     {rob_uop_19_uses_stq},
     {rob_uop_18_uses_stq},
     {rob_uop_17_uses_stq},
     {rob_uop_16_uses_stq},
     {rob_uop_15_uses_stq},
     {rob_uop_14_uses_stq},
     {rob_uop_13_uses_stq},
     {rob_uop_12_uses_stq},
     {rob_uop_11_uses_stq},
     {rob_uop_10_uses_stq},
     {rob_uop_9_uses_stq},
     {rob_uop_8_uses_stq},
     {rob_uop_7_uses_stq},
     {rob_uop_6_uses_stq},
     {rob_uop_5_uses_stq},
     {rob_uop_4_uses_stq},
     {rob_uop_3_uses_stq},
     {rob_uop_2_uses_stq},
     {rob_uop_1_uses_stq},
     {rob_uop_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_23 =
    {{rob_uop_31_is_sys_pc2epc},
     {rob_uop_30_is_sys_pc2epc},
     {rob_uop_29_is_sys_pc2epc},
     {rob_uop_28_is_sys_pc2epc},
     {rob_uop_27_is_sys_pc2epc},
     {rob_uop_26_is_sys_pc2epc},
     {rob_uop_25_is_sys_pc2epc},
     {rob_uop_24_is_sys_pc2epc},
     {rob_uop_23_is_sys_pc2epc},
     {rob_uop_22_is_sys_pc2epc},
     {rob_uop_21_is_sys_pc2epc},
     {rob_uop_20_is_sys_pc2epc},
     {rob_uop_19_is_sys_pc2epc},
     {rob_uop_18_is_sys_pc2epc},
     {rob_uop_17_is_sys_pc2epc},
     {rob_uop_16_is_sys_pc2epc},
     {rob_uop_15_is_sys_pc2epc},
     {rob_uop_14_is_sys_pc2epc},
     {rob_uop_13_is_sys_pc2epc},
     {rob_uop_12_is_sys_pc2epc},
     {rob_uop_11_is_sys_pc2epc},
     {rob_uop_10_is_sys_pc2epc},
     {rob_uop_9_is_sys_pc2epc},
     {rob_uop_8_is_sys_pc2epc},
     {rob_uop_7_is_sys_pc2epc},
     {rob_uop_6_is_sys_pc2epc},
     {rob_uop_5_is_sys_pc2epc},
     {rob_uop_4_is_sys_pc2epc},
     {rob_uop_3_is_sys_pc2epc},
     {rob_uop_2_is_sys_pc2epc},
     {rob_uop_1_is_sys_pc2epc},
     {rob_uop_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_24 =
    {{rob_uop_31_flush_on_commit},
     {rob_uop_30_flush_on_commit},
     {rob_uop_29_flush_on_commit},
     {rob_uop_28_flush_on_commit},
     {rob_uop_27_flush_on_commit},
     {rob_uop_26_flush_on_commit},
     {rob_uop_25_flush_on_commit},
     {rob_uop_24_flush_on_commit},
     {rob_uop_23_flush_on_commit},
     {rob_uop_22_flush_on_commit},
     {rob_uop_21_flush_on_commit},
     {rob_uop_20_flush_on_commit},
     {rob_uop_19_flush_on_commit},
     {rob_uop_18_flush_on_commit},
     {rob_uop_17_flush_on_commit},
     {rob_uop_16_flush_on_commit},
     {rob_uop_15_flush_on_commit},
     {rob_uop_14_flush_on_commit},
     {rob_uop_13_flush_on_commit},
     {rob_uop_12_flush_on_commit},
     {rob_uop_11_flush_on_commit},
     {rob_uop_10_flush_on_commit},
     {rob_uop_9_flush_on_commit},
     {rob_uop_8_flush_on_commit},
     {rob_uop_7_flush_on_commit},
     {rob_uop_6_flush_on_commit},
     {rob_uop_5_flush_on_commit},
     {rob_uop_4_flush_on_commit},
     {rob_uop_3_flush_on_commit},
     {rob_uop_2_flush_on_commit},
     {rob_uop_1_flush_on_commit},
     {rob_uop_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_25 =
    {{rob_uop_31_ldst},
     {rob_uop_30_ldst},
     {rob_uop_29_ldst},
     {rob_uop_28_ldst},
     {rob_uop_27_ldst},
     {rob_uop_26_ldst},
     {rob_uop_25_ldst},
     {rob_uop_24_ldst},
     {rob_uop_23_ldst},
     {rob_uop_22_ldst},
     {rob_uop_21_ldst},
     {rob_uop_20_ldst},
     {rob_uop_19_ldst},
     {rob_uop_18_ldst},
     {rob_uop_17_ldst},
     {rob_uop_16_ldst},
     {rob_uop_15_ldst},
     {rob_uop_14_ldst},
     {rob_uop_13_ldst},
     {rob_uop_12_ldst},
     {rob_uop_11_ldst},
     {rob_uop_10_ldst},
     {rob_uop_9_ldst},
     {rob_uop_8_ldst},
     {rob_uop_7_ldst},
     {rob_uop_6_ldst},
     {rob_uop_5_ldst},
     {rob_uop_4_ldst},
     {rob_uop_3_ldst},
     {rob_uop_2_ldst},
     {rob_uop_1_ldst},
     {rob_uop_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_26 =
    {{rob_uop_31_ldst_val},
     {rob_uop_30_ldst_val},
     {rob_uop_29_ldst_val},
     {rob_uop_28_ldst_val},
     {rob_uop_27_ldst_val},
     {rob_uop_26_ldst_val},
     {rob_uop_25_ldst_val},
     {rob_uop_24_ldst_val},
     {rob_uop_23_ldst_val},
     {rob_uop_22_ldst_val},
     {rob_uop_21_ldst_val},
     {rob_uop_20_ldst_val},
     {rob_uop_19_ldst_val},
     {rob_uop_18_ldst_val},
     {rob_uop_17_ldst_val},
     {rob_uop_16_ldst_val},
     {rob_uop_15_ldst_val},
     {rob_uop_14_ldst_val},
     {rob_uop_13_ldst_val},
     {rob_uop_12_ldst_val},
     {rob_uop_11_ldst_val},
     {rob_uop_10_ldst_val},
     {rob_uop_9_ldst_val},
     {rob_uop_8_ldst_val},
     {rob_uop_7_ldst_val},
     {rob_uop_6_ldst_val},
     {rob_uop_5_ldst_val},
     {rob_uop_4_ldst_val},
     {rob_uop_3_ldst_val},
     {rob_uop_2_ldst_val},
     {rob_uop_1_ldst_val},
     {rob_uop_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_27 =
    {{rob_uop_31_dst_rtype},
     {rob_uop_30_dst_rtype},
     {rob_uop_29_dst_rtype},
     {rob_uop_28_dst_rtype},
     {rob_uop_27_dst_rtype},
     {rob_uop_26_dst_rtype},
     {rob_uop_25_dst_rtype},
     {rob_uop_24_dst_rtype},
     {rob_uop_23_dst_rtype},
     {rob_uop_22_dst_rtype},
     {rob_uop_21_dst_rtype},
     {rob_uop_20_dst_rtype},
     {rob_uop_19_dst_rtype},
     {rob_uop_18_dst_rtype},
     {rob_uop_17_dst_rtype},
     {rob_uop_16_dst_rtype},
     {rob_uop_15_dst_rtype},
     {rob_uop_14_dst_rtype},
     {rob_uop_13_dst_rtype},
     {rob_uop_12_dst_rtype},
     {rob_uop_11_dst_rtype},
     {rob_uop_10_dst_rtype},
     {rob_uop_9_dst_rtype},
     {rob_uop_8_dst_rtype},
     {rob_uop_7_dst_rtype},
     {rob_uop_6_dst_rtype},
     {rob_uop_5_dst_rtype},
     {rob_uop_4_dst_rtype},
     {rob_uop_3_dst_rtype},
     {rob_uop_2_dst_rtype},
     {rob_uop_1_dst_rtype},
     {rob_uop_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_28 =
    {{rob_uop_31_fp_val},
     {rob_uop_30_fp_val},
     {rob_uop_29_fp_val},
     {rob_uop_28_fp_val},
     {rob_uop_27_fp_val},
     {rob_uop_26_fp_val},
     {rob_uop_25_fp_val},
     {rob_uop_24_fp_val},
     {rob_uop_23_fp_val},
     {rob_uop_22_fp_val},
     {rob_uop_21_fp_val},
     {rob_uop_20_fp_val},
     {rob_uop_19_fp_val},
     {rob_uop_18_fp_val},
     {rob_uop_17_fp_val},
     {rob_uop_16_fp_val},
     {rob_uop_15_fp_val},
     {rob_uop_14_fp_val},
     {rob_uop_13_fp_val},
     {rob_uop_12_fp_val},
     {rob_uop_11_fp_val},
     {rob_uop_10_fp_val},
     {rob_uop_9_fp_val},
     {rob_uop_8_fp_val},
     {rob_uop_7_fp_val},
     {rob_uop_6_fp_val},
     {rob_uop_5_fp_val},
     {rob_uop_4_fp_val},
     {rob_uop_3_fp_val},
     {rob_uop_2_fp_val},
     {rob_uop_1_fp_val},
     {rob_uop_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row = _io_commit_rollback_T_2 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_0_output = rbk_row & _GEN[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              rob_val_1_0;	// rob.scala:307:32
  reg              rob_val_1_1;	// rob.scala:307:32
  reg              rob_val_1_2;	// rob.scala:307:32
  reg              rob_val_1_3;	// rob.scala:307:32
  reg              rob_val_1_4;	// rob.scala:307:32
  reg              rob_val_1_5;	// rob.scala:307:32
  reg              rob_val_1_6;	// rob.scala:307:32
  reg              rob_val_1_7;	// rob.scala:307:32
  reg              rob_val_1_8;	// rob.scala:307:32
  reg              rob_val_1_9;	// rob.scala:307:32
  reg              rob_val_1_10;	// rob.scala:307:32
  reg              rob_val_1_11;	// rob.scala:307:32
  reg              rob_val_1_12;	// rob.scala:307:32
  reg              rob_val_1_13;	// rob.scala:307:32
  reg              rob_val_1_14;	// rob.scala:307:32
  reg              rob_val_1_15;	// rob.scala:307:32
  reg              rob_val_1_16;	// rob.scala:307:32
  reg              rob_val_1_17;	// rob.scala:307:32
  reg              rob_val_1_18;	// rob.scala:307:32
  reg              rob_val_1_19;	// rob.scala:307:32
  reg              rob_val_1_20;	// rob.scala:307:32
  reg              rob_val_1_21;	// rob.scala:307:32
  reg              rob_val_1_22;	// rob.scala:307:32
  reg              rob_val_1_23;	// rob.scala:307:32
  reg              rob_val_1_24;	// rob.scala:307:32
  reg              rob_val_1_25;	// rob.scala:307:32
  reg              rob_val_1_26;	// rob.scala:307:32
  reg              rob_val_1_27;	// rob.scala:307:32
  reg              rob_val_1_28;	// rob.scala:307:32
  reg              rob_val_1_29;	// rob.scala:307:32
  reg              rob_val_1_30;	// rob.scala:307:32
  reg              rob_val_1_31;	// rob.scala:307:32
  reg              rob_bsy_1_0;	// rob.scala:308:28
  reg              rob_bsy_1_1;	// rob.scala:308:28
  reg              rob_bsy_1_2;	// rob.scala:308:28
  reg              rob_bsy_1_3;	// rob.scala:308:28
  reg              rob_bsy_1_4;	// rob.scala:308:28
  reg              rob_bsy_1_5;	// rob.scala:308:28
  reg              rob_bsy_1_6;	// rob.scala:308:28
  reg              rob_bsy_1_7;	// rob.scala:308:28
  reg              rob_bsy_1_8;	// rob.scala:308:28
  reg              rob_bsy_1_9;	// rob.scala:308:28
  reg              rob_bsy_1_10;	// rob.scala:308:28
  reg              rob_bsy_1_11;	// rob.scala:308:28
  reg              rob_bsy_1_12;	// rob.scala:308:28
  reg              rob_bsy_1_13;	// rob.scala:308:28
  reg              rob_bsy_1_14;	// rob.scala:308:28
  reg              rob_bsy_1_15;	// rob.scala:308:28
  reg              rob_bsy_1_16;	// rob.scala:308:28
  reg              rob_bsy_1_17;	// rob.scala:308:28
  reg              rob_bsy_1_18;	// rob.scala:308:28
  reg              rob_bsy_1_19;	// rob.scala:308:28
  reg              rob_bsy_1_20;	// rob.scala:308:28
  reg              rob_bsy_1_21;	// rob.scala:308:28
  reg              rob_bsy_1_22;	// rob.scala:308:28
  reg              rob_bsy_1_23;	// rob.scala:308:28
  reg              rob_bsy_1_24;	// rob.scala:308:28
  reg              rob_bsy_1_25;	// rob.scala:308:28
  reg              rob_bsy_1_26;	// rob.scala:308:28
  reg              rob_bsy_1_27;	// rob.scala:308:28
  reg              rob_bsy_1_28;	// rob.scala:308:28
  reg              rob_bsy_1_29;	// rob.scala:308:28
  reg              rob_bsy_1_30;	// rob.scala:308:28
  reg              rob_bsy_1_31;	// rob.scala:308:28
  reg              rob_unsafe_1_0;	// rob.scala:309:28
  reg              rob_unsafe_1_1;	// rob.scala:309:28
  reg              rob_unsafe_1_2;	// rob.scala:309:28
  reg              rob_unsafe_1_3;	// rob.scala:309:28
  reg              rob_unsafe_1_4;	// rob.scala:309:28
  reg              rob_unsafe_1_5;	// rob.scala:309:28
  reg              rob_unsafe_1_6;	// rob.scala:309:28
  reg              rob_unsafe_1_7;	// rob.scala:309:28
  reg              rob_unsafe_1_8;	// rob.scala:309:28
  reg              rob_unsafe_1_9;	// rob.scala:309:28
  reg              rob_unsafe_1_10;	// rob.scala:309:28
  reg              rob_unsafe_1_11;	// rob.scala:309:28
  reg              rob_unsafe_1_12;	// rob.scala:309:28
  reg              rob_unsafe_1_13;	// rob.scala:309:28
  reg              rob_unsafe_1_14;	// rob.scala:309:28
  reg              rob_unsafe_1_15;	// rob.scala:309:28
  reg              rob_unsafe_1_16;	// rob.scala:309:28
  reg              rob_unsafe_1_17;	// rob.scala:309:28
  reg              rob_unsafe_1_18;	// rob.scala:309:28
  reg              rob_unsafe_1_19;	// rob.scala:309:28
  reg              rob_unsafe_1_20;	// rob.scala:309:28
  reg              rob_unsafe_1_21;	// rob.scala:309:28
  reg              rob_unsafe_1_22;	// rob.scala:309:28
  reg              rob_unsafe_1_23;	// rob.scala:309:28
  reg              rob_unsafe_1_24;	// rob.scala:309:28
  reg              rob_unsafe_1_25;	// rob.scala:309:28
  reg              rob_unsafe_1_26;	// rob.scala:309:28
  reg              rob_unsafe_1_27;	// rob.scala:309:28
  reg              rob_unsafe_1_28;	// rob.scala:309:28
  reg              rob_unsafe_1_29;	// rob.scala:309:28
  reg              rob_unsafe_1_30;	// rob.scala:309:28
  reg              rob_unsafe_1_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_1_0_uopc;	// rob.scala:310:28
  reg              rob_uop_1_0_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_0_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_0_ldst;	// rob.scala:310:28
  reg              rob_uop_1_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_1_uopc;	// rob.scala:310:28
  reg              rob_uop_1_1_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_1_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_1_ldst;	// rob.scala:310:28
  reg              rob_uop_1_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_2_uopc;	// rob.scala:310:28
  reg              rob_uop_1_2_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_2_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_2_ldst;	// rob.scala:310:28
  reg              rob_uop_1_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_3_uopc;	// rob.scala:310:28
  reg              rob_uop_1_3_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_3_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_3_ldst;	// rob.scala:310:28
  reg              rob_uop_1_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_4_uopc;	// rob.scala:310:28
  reg              rob_uop_1_4_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_4_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_4_ldst;	// rob.scala:310:28
  reg              rob_uop_1_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_5_uopc;	// rob.scala:310:28
  reg              rob_uop_1_5_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_5_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_5_ldst;	// rob.scala:310:28
  reg              rob_uop_1_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_6_uopc;	// rob.scala:310:28
  reg              rob_uop_1_6_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_6_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_6_ldst;	// rob.scala:310:28
  reg              rob_uop_1_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_7_uopc;	// rob.scala:310:28
  reg              rob_uop_1_7_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_7_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_7_ldst;	// rob.scala:310:28
  reg              rob_uop_1_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_8_uopc;	// rob.scala:310:28
  reg              rob_uop_1_8_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_8_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_8_ldst;	// rob.scala:310:28
  reg              rob_uop_1_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_9_uopc;	// rob.scala:310:28
  reg              rob_uop_1_9_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_9_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_9_ldst;	// rob.scala:310:28
  reg              rob_uop_1_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_10_uopc;	// rob.scala:310:28
  reg              rob_uop_1_10_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_10_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_10_ldst;	// rob.scala:310:28
  reg              rob_uop_1_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_11_uopc;	// rob.scala:310:28
  reg              rob_uop_1_11_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_11_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_11_ldst;	// rob.scala:310:28
  reg              rob_uop_1_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_12_uopc;	// rob.scala:310:28
  reg              rob_uop_1_12_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_12_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_12_ldst;	// rob.scala:310:28
  reg              rob_uop_1_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_13_uopc;	// rob.scala:310:28
  reg              rob_uop_1_13_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_13_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_13_ldst;	// rob.scala:310:28
  reg              rob_uop_1_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_14_uopc;	// rob.scala:310:28
  reg              rob_uop_1_14_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_14_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_14_ldst;	// rob.scala:310:28
  reg              rob_uop_1_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_15_uopc;	// rob.scala:310:28
  reg              rob_uop_1_15_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_15_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_15_ldst;	// rob.scala:310:28
  reg              rob_uop_1_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_16_uopc;	// rob.scala:310:28
  reg              rob_uop_1_16_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_16_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_16_ldst;	// rob.scala:310:28
  reg              rob_uop_1_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_17_uopc;	// rob.scala:310:28
  reg              rob_uop_1_17_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_17_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_17_ldst;	// rob.scala:310:28
  reg              rob_uop_1_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_18_uopc;	// rob.scala:310:28
  reg              rob_uop_1_18_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_18_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_18_ldst;	// rob.scala:310:28
  reg              rob_uop_1_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_19_uopc;	// rob.scala:310:28
  reg              rob_uop_1_19_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_19_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_19_ldst;	// rob.scala:310:28
  reg              rob_uop_1_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_20_uopc;	// rob.scala:310:28
  reg              rob_uop_1_20_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_20_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_20_ldst;	// rob.scala:310:28
  reg              rob_uop_1_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_21_uopc;	// rob.scala:310:28
  reg              rob_uop_1_21_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_21_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_21_ldst;	// rob.scala:310:28
  reg              rob_uop_1_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_22_uopc;	// rob.scala:310:28
  reg              rob_uop_1_22_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_22_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_22_ldst;	// rob.scala:310:28
  reg              rob_uop_1_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_23_uopc;	// rob.scala:310:28
  reg              rob_uop_1_23_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_23_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_23_ldst;	// rob.scala:310:28
  reg              rob_uop_1_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_24_uopc;	// rob.scala:310:28
  reg              rob_uop_1_24_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_24_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_24_ldst;	// rob.scala:310:28
  reg              rob_uop_1_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_25_uopc;	// rob.scala:310:28
  reg              rob_uop_1_25_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_25_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_25_ldst;	// rob.scala:310:28
  reg              rob_uop_1_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_26_uopc;	// rob.scala:310:28
  reg              rob_uop_1_26_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_26_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_26_ldst;	// rob.scala:310:28
  reg              rob_uop_1_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_27_uopc;	// rob.scala:310:28
  reg              rob_uop_1_27_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_27_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_27_ldst;	// rob.scala:310:28
  reg              rob_uop_1_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_28_uopc;	// rob.scala:310:28
  reg              rob_uop_1_28_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_28_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_28_ldst;	// rob.scala:310:28
  reg              rob_uop_1_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_29_uopc;	// rob.scala:310:28
  reg              rob_uop_1_29_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_29_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_29_ldst;	// rob.scala:310:28
  reg              rob_uop_1_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_30_uopc;	// rob.scala:310:28
  reg              rob_uop_1_30_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_30_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_30_ldst;	// rob.scala:310:28
  reg              rob_uop_1_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_31_uopc;	// rob.scala:310:28
  reg              rob_uop_1_31_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_1_31_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_1_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_1_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_1_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_1_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_1_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_1_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_1_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_1_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_1_31_ldst;	// rob.scala:310:28
  reg              rob_uop_1_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_1_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_1_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_1_0;	// rob.scala:311:28
  reg              rob_exception_1_1;	// rob.scala:311:28
  reg              rob_exception_1_2;	// rob.scala:311:28
  reg              rob_exception_1_3;	// rob.scala:311:28
  reg              rob_exception_1_4;	// rob.scala:311:28
  reg              rob_exception_1_5;	// rob.scala:311:28
  reg              rob_exception_1_6;	// rob.scala:311:28
  reg              rob_exception_1_7;	// rob.scala:311:28
  reg              rob_exception_1_8;	// rob.scala:311:28
  reg              rob_exception_1_9;	// rob.scala:311:28
  reg              rob_exception_1_10;	// rob.scala:311:28
  reg              rob_exception_1_11;	// rob.scala:311:28
  reg              rob_exception_1_12;	// rob.scala:311:28
  reg              rob_exception_1_13;	// rob.scala:311:28
  reg              rob_exception_1_14;	// rob.scala:311:28
  reg              rob_exception_1_15;	// rob.scala:311:28
  reg              rob_exception_1_16;	// rob.scala:311:28
  reg              rob_exception_1_17;	// rob.scala:311:28
  reg              rob_exception_1_18;	// rob.scala:311:28
  reg              rob_exception_1_19;	// rob.scala:311:28
  reg              rob_exception_1_20;	// rob.scala:311:28
  reg              rob_exception_1_21;	// rob.scala:311:28
  reg              rob_exception_1_22;	// rob.scala:311:28
  reg              rob_exception_1_23;	// rob.scala:311:28
  reg              rob_exception_1_24;	// rob.scala:311:28
  reg              rob_exception_1_25;	// rob.scala:311:28
  reg              rob_exception_1_26;	// rob.scala:311:28
  reg              rob_exception_1_27;	// rob.scala:311:28
  reg              rob_exception_1_28;	// rob.scala:311:28
  reg              rob_exception_1_29;	// rob.scala:311:28
  reg              rob_exception_1_30;	// rob.scala:311:28
  reg              rob_exception_1_31;	// rob.scala:311:28
  reg              rob_predicated_1_0;	// rob.scala:312:29
  reg              rob_predicated_1_1;	// rob.scala:312:29
  reg              rob_predicated_1_2;	// rob.scala:312:29
  reg              rob_predicated_1_3;	// rob.scala:312:29
  reg              rob_predicated_1_4;	// rob.scala:312:29
  reg              rob_predicated_1_5;	// rob.scala:312:29
  reg              rob_predicated_1_6;	// rob.scala:312:29
  reg              rob_predicated_1_7;	// rob.scala:312:29
  reg              rob_predicated_1_8;	// rob.scala:312:29
  reg              rob_predicated_1_9;	// rob.scala:312:29
  reg              rob_predicated_1_10;	// rob.scala:312:29
  reg              rob_predicated_1_11;	// rob.scala:312:29
  reg              rob_predicated_1_12;	// rob.scala:312:29
  reg              rob_predicated_1_13;	// rob.scala:312:29
  reg              rob_predicated_1_14;	// rob.scala:312:29
  reg              rob_predicated_1_15;	// rob.scala:312:29
  reg              rob_predicated_1_16;	// rob.scala:312:29
  reg              rob_predicated_1_17;	// rob.scala:312:29
  reg              rob_predicated_1_18;	// rob.scala:312:29
  reg              rob_predicated_1_19;	// rob.scala:312:29
  reg              rob_predicated_1_20;	// rob.scala:312:29
  reg              rob_predicated_1_21;	// rob.scala:312:29
  reg              rob_predicated_1_22;	// rob.scala:312:29
  reg              rob_predicated_1_23;	// rob.scala:312:29
  reg              rob_predicated_1_24;	// rob.scala:312:29
  reg              rob_predicated_1_25;	// rob.scala:312:29
  reg              rob_predicated_1_26;	// rob.scala:312:29
  reg              rob_predicated_1_27;	// rob.scala:312:29
  reg              rob_predicated_1_28;	// rob.scala:312:29
  reg              rob_predicated_1_29;	// rob.scala:312:29
  reg              rob_predicated_1_30;	// rob.scala:312:29
  reg              rob_predicated_1_31;	// rob.scala:312:29
  wire [31:0]      _GEN_29 =
    {{rob_val_1_31},
     {rob_val_1_30},
     {rob_val_1_29},
     {rob_val_1_28},
     {rob_val_1_27},
     {rob_val_1_26},
     {rob_val_1_25},
     {rob_val_1_24},
     {rob_val_1_23},
     {rob_val_1_22},
     {rob_val_1_21},
     {rob_val_1_20},
     {rob_val_1_19},
     {rob_val_1_18},
     {rob_val_1_17},
     {rob_val_1_16},
     {rob_val_1_15},
     {rob_val_1_14},
     {rob_val_1_13},
     {rob_val_1_12},
     {rob_val_1_11},
     {rob_val_1_10},
     {rob_val_1_9},
     {rob_val_1_8},
     {rob_val_1_7},
     {rob_val_1_6},
     {rob_val_1_5},
     {rob_val_1_4},
     {rob_val_1_3},
     {rob_val_1_2},
     {rob_val_1_1},
     {rob_val_1_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_1 = _GEN_29[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_30 =
    io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_31 =
    io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_32 =
    io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_33 =
    io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_34 =
    io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_35 =
    io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :346:27, :540:33
  wire             _GEN_36 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :361:31, :540:33
  wire [31:0]      _GEN_37 =
    {{rob_bsy_1_31},
     {rob_bsy_1_30},
     {rob_bsy_1_29},
     {rob_bsy_1_28},
     {rob_bsy_1_27},
     {rob_bsy_1_26},
     {rob_bsy_1_25},
     {rob_bsy_1_24},
     {rob_bsy_1_23},
     {rob_bsy_1_22},
     {rob_bsy_1_21},
     {rob_bsy_1_20},
     {rob_bsy_1_19},
     {rob_bsy_1_18},
     {rob_bsy_1_17},
     {rob_bsy_1_16},
     {rob_bsy_1_15},
     {rob_bsy_1_14},
     {rob_bsy_1_13},
     {rob_bsy_1_12},
     {rob_bsy_1_11},
     {rob_bsy_1_10},
     {rob_bsy_1_9},
     {rob_bsy_1_8},
     {rob_bsy_1_7},
     {rob_bsy_1_6},
     {rob_bsy_1_5},
     {rob_bsy_1_4},
     {rob_bsy_1_3},
     {rob_bsy_1_2},
     {rob_bsy_1_1},
     {rob_bsy_1_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_38 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :361:31, :540:33
  wire             _GEN_39 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h1;	// rob.scala:272:36, :304:53, :390:26, :540:33
  wire [31:0]      _GEN_40 =
    {{rob_unsafe_1_31},
     {rob_unsafe_1_30},
     {rob_unsafe_1_29},
     {rob_unsafe_1_28},
     {rob_unsafe_1_27},
     {rob_unsafe_1_26},
     {rob_unsafe_1_25},
     {rob_unsafe_1_24},
     {rob_unsafe_1_23},
     {rob_unsafe_1_22},
     {rob_unsafe_1_21},
     {rob_unsafe_1_20},
     {rob_unsafe_1_19},
     {rob_unsafe_1_18},
     {rob_unsafe_1_17},
     {rob_unsafe_1_16},
     {rob_unsafe_1_15},
     {rob_unsafe_1_14},
     {rob_unsafe_1_13},
     {rob_unsafe_1_12},
     {rob_unsafe_1_11},
     {rob_unsafe_1_10},
     {rob_unsafe_1_9},
     {rob_unsafe_1_8},
     {rob_unsafe_1_7},
     {rob_unsafe_1_6},
     {rob_unsafe_1_5},
     {rob_unsafe_1_4},
     {rob_unsafe_1_3},
     {rob_unsafe_1_2},
     {rob_unsafe_1_1},
     {rob_unsafe_1_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_1 = _GEN_29[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_41 =
    {{rob_exception_1_31},
     {rob_exception_1_30},
     {rob_exception_1_29},
     {rob_exception_1_28},
     {rob_exception_1_27},
     {rob_exception_1_26},
     {rob_exception_1_25},
     {rob_exception_1_24},
     {rob_exception_1_23},
     {rob_exception_1_22},
     {rob_exception_1_21},
     {rob_exception_1_20},
     {rob_exception_1_19},
     {rob_exception_1_18},
     {rob_exception_1_17},
     {rob_exception_1_16},
     {rob_exception_1_15},
     {rob_exception_1_14},
     {rob_exception_1_13},
     {rob_exception_1_12},
     {rob_exception_1_11},
     {rob_exception_1_10},
     {rob_exception_1_9},
     {rob_exception_1_8},
     {rob_exception_1_7},
     {rob_exception_1_6},
     {rob_exception_1_5},
     {rob_exception_1_4},
     {rob_exception_1_3},
     {rob_exception_1_2},
     {rob_exception_1_1},
     {rob_exception_1_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_1 = rob_head_vals_1 & _GEN_41[rob_head];	// rob.scala:224:29, :398:49
  wire             can_commit_1 = rob_head_vals_1 & ~_GEN_37[rob_head] & ~io_csr_stall;	// rob.scala:224:29, :366:31, :398:49, :404:{43,64,67}
  wire [31:0]      _GEN_42 =
    {{rob_predicated_1_31},
     {rob_predicated_1_30},
     {rob_predicated_1_29},
     {rob_predicated_1_28},
     {rob_predicated_1_27},
     {rob_predicated_1_26},
     {rob_predicated_1_25},
     {rob_predicated_1_24},
     {rob_predicated_1_23},
     {rob_predicated_1_22},
     {rob_predicated_1_21},
     {rob_predicated_1_20},
     {rob_predicated_1_19},
     {rob_predicated_1_18},
     {rob_predicated_1_17},
     {rob_predicated_1_16},
     {rob_predicated_1_15},
     {rob_predicated_1_14},
     {rob_predicated_1_13},
     {rob_predicated_1_12},
     {rob_predicated_1_11},
     {rob_predicated_1_10},
     {rob_predicated_1_9},
     {rob_predicated_1_8},
     {rob_predicated_1_7},
     {rob_predicated_1_6},
     {rob_predicated_1_5},
     {rob_predicated_1_4},
     {rob_predicated_1_3},
     {rob_predicated_1_2},
     {rob_predicated_1_1},
     {rob_predicated_1_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_43 =
    {{rob_uop_1_31_uopc},
     {rob_uop_1_30_uopc},
     {rob_uop_1_29_uopc},
     {rob_uop_1_28_uopc},
     {rob_uop_1_27_uopc},
     {rob_uop_1_26_uopc},
     {rob_uop_1_25_uopc},
     {rob_uop_1_24_uopc},
     {rob_uop_1_23_uopc},
     {rob_uop_1_22_uopc},
     {rob_uop_1_21_uopc},
     {rob_uop_1_20_uopc},
     {rob_uop_1_19_uopc},
     {rob_uop_1_18_uopc},
     {rob_uop_1_17_uopc},
     {rob_uop_1_16_uopc},
     {rob_uop_1_15_uopc},
     {rob_uop_1_14_uopc},
     {rob_uop_1_13_uopc},
     {rob_uop_1_12_uopc},
     {rob_uop_1_11_uopc},
     {rob_uop_1_10_uopc},
     {rob_uop_1_9_uopc},
     {rob_uop_1_8_uopc},
     {rob_uop_1_7_uopc},
     {rob_uop_1_6_uopc},
     {rob_uop_1_5_uopc},
     {rob_uop_1_4_uopc},
     {rob_uop_1_3_uopc},
     {rob_uop_1_2_uopc},
     {rob_uop_1_1_uopc},
     {rob_uop_1_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_44 =
    {{rob_uop_1_31_is_rvc},
     {rob_uop_1_30_is_rvc},
     {rob_uop_1_29_is_rvc},
     {rob_uop_1_28_is_rvc},
     {rob_uop_1_27_is_rvc},
     {rob_uop_1_26_is_rvc},
     {rob_uop_1_25_is_rvc},
     {rob_uop_1_24_is_rvc},
     {rob_uop_1_23_is_rvc},
     {rob_uop_1_22_is_rvc},
     {rob_uop_1_21_is_rvc},
     {rob_uop_1_20_is_rvc},
     {rob_uop_1_19_is_rvc},
     {rob_uop_1_18_is_rvc},
     {rob_uop_1_17_is_rvc},
     {rob_uop_1_16_is_rvc},
     {rob_uop_1_15_is_rvc},
     {rob_uop_1_14_is_rvc},
     {rob_uop_1_13_is_rvc},
     {rob_uop_1_12_is_rvc},
     {rob_uop_1_11_is_rvc},
     {rob_uop_1_10_is_rvc},
     {rob_uop_1_9_is_rvc},
     {rob_uop_1_8_is_rvc},
     {rob_uop_1_7_is_rvc},
     {rob_uop_1_6_is_rvc},
     {rob_uop_1_5_is_rvc},
     {rob_uop_1_4_is_rvc},
     {rob_uop_1_3_is_rvc},
     {rob_uop_1_2_is_rvc},
     {rob_uop_1_1_is_rvc},
     {rob_uop_1_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][4:0] _GEN_45 =
    {{rob_uop_1_31_ftq_idx},
     {rob_uop_1_30_ftq_idx},
     {rob_uop_1_29_ftq_idx},
     {rob_uop_1_28_ftq_idx},
     {rob_uop_1_27_ftq_idx},
     {rob_uop_1_26_ftq_idx},
     {rob_uop_1_25_ftq_idx},
     {rob_uop_1_24_ftq_idx},
     {rob_uop_1_23_ftq_idx},
     {rob_uop_1_22_ftq_idx},
     {rob_uop_1_21_ftq_idx},
     {rob_uop_1_20_ftq_idx},
     {rob_uop_1_19_ftq_idx},
     {rob_uop_1_18_ftq_idx},
     {rob_uop_1_17_ftq_idx},
     {rob_uop_1_16_ftq_idx},
     {rob_uop_1_15_ftq_idx},
     {rob_uop_1_14_ftq_idx},
     {rob_uop_1_13_ftq_idx},
     {rob_uop_1_12_ftq_idx},
     {rob_uop_1_11_ftq_idx},
     {rob_uop_1_10_ftq_idx},
     {rob_uop_1_9_ftq_idx},
     {rob_uop_1_8_ftq_idx},
     {rob_uop_1_7_ftq_idx},
     {rob_uop_1_6_ftq_idx},
     {rob_uop_1_5_ftq_idx},
     {rob_uop_1_4_ftq_idx},
     {rob_uop_1_3_ftq_idx},
     {rob_uop_1_2_ftq_idx},
     {rob_uop_1_1_ftq_idx},
     {rob_uop_1_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_46 =
    {{rob_uop_1_31_edge_inst},
     {rob_uop_1_30_edge_inst},
     {rob_uop_1_29_edge_inst},
     {rob_uop_1_28_edge_inst},
     {rob_uop_1_27_edge_inst},
     {rob_uop_1_26_edge_inst},
     {rob_uop_1_25_edge_inst},
     {rob_uop_1_24_edge_inst},
     {rob_uop_1_23_edge_inst},
     {rob_uop_1_22_edge_inst},
     {rob_uop_1_21_edge_inst},
     {rob_uop_1_20_edge_inst},
     {rob_uop_1_19_edge_inst},
     {rob_uop_1_18_edge_inst},
     {rob_uop_1_17_edge_inst},
     {rob_uop_1_16_edge_inst},
     {rob_uop_1_15_edge_inst},
     {rob_uop_1_14_edge_inst},
     {rob_uop_1_13_edge_inst},
     {rob_uop_1_12_edge_inst},
     {rob_uop_1_11_edge_inst},
     {rob_uop_1_10_edge_inst},
     {rob_uop_1_9_edge_inst},
     {rob_uop_1_8_edge_inst},
     {rob_uop_1_7_edge_inst},
     {rob_uop_1_6_edge_inst},
     {rob_uop_1_5_edge_inst},
     {rob_uop_1_4_edge_inst},
     {rob_uop_1_3_edge_inst},
     {rob_uop_1_2_edge_inst},
     {rob_uop_1_1_edge_inst},
     {rob_uop_1_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_47 =
    {{rob_uop_1_31_pc_lob},
     {rob_uop_1_30_pc_lob},
     {rob_uop_1_29_pc_lob},
     {rob_uop_1_28_pc_lob},
     {rob_uop_1_27_pc_lob},
     {rob_uop_1_26_pc_lob},
     {rob_uop_1_25_pc_lob},
     {rob_uop_1_24_pc_lob},
     {rob_uop_1_23_pc_lob},
     {rob_uop_1_22_pc_lob},
     {rob_uop_1_21_pc_lob},
     {rob_uop_1_20_pc_lob},
     {rob_uop_1_19_pc_lob},
     {rob_uop_1_18_pc_lob},
     {rob_uop_1_17_pc_lob},
     {rob_uop_1_16_pc_lob},
     {rob_uop_1_15_pc_lob},
     {rob_uop_1_14_pc_lob},
     {rob_uop_1_13_pc_lob},
     {rob_uop_1_12_pc_lob},
     {rob_uop_1_11_pc_lob},
     {rob_uop_1_10_pc_lob},
     {rob_uop_1_9_pc_lob},
     {rob_uop_1_8_pc_lob},
     {rob_uop_1_7_pc_lob},
     {rob_uop_1_6_pc_lob},
     {rob_uop_1_5_pc_lob},
     {rob_uop_1_4_pc_lob},
     {rob_uop_1_3_pc_lob},
     {rob_uop_1_2_pc_lob},
     {rob_uop_1_1_pc_lob},
     {rob_uop_1_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_48 =
    {{rob_uop_1_31_pdst},
     {rob_uop_1_30_pdst},
     {rob_uop_1_29_pdst},
     {rob_uop_1_28_pdst},
     {rob_uop_1_27_pdst},
     {rob_uop_1_26_pdst},
     {rob_uop_1_25_pdst},
     {rob_uop_1_24_pdst},
     {rob_uop_1_23_pdst},
     {rob_uop_1_22_pdst},
     {rob_uop_1_21_pdst},
     {rob_uop_1_20_pdst},
     {rob_uop_1_19_pdst},
     {rob_uop_1_18_pdst},
     {rob_uop_1_17_pdst},
     {rob_uop_1_16_pdst},
     {rob_uop_1_15_pdst},
     {rob_uop_1_14_pdst},
     {rob_uop_1_13_pdst},
     {rob_uop_1_12_pdst},
     {rob_uop_1_11_pdst},
     {rob_uop_1_10_pdst},
     {rob_uop_1_9_pdst},
     {rob_uop_1_8_pdst},
     {rob_uop_1_7_pdst},
     {rob_uop_1_6_pdst},
     {rob_uop_1_5_pdst},
     {rob_uop_1_4_pdst},
     {rob_uop_1_3_pdst},
     {rob_uop_1_2_pdst},
     {rob_uop_1_1_pdst},
     {rob_uop_1_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_49 =
    {{rob_uop_1_31_stale_pdst},
     {rob_uop_1_30_stale_pdst},
     {rob_uop_1_29_stale_pdst},
     {rob_uop_1_28_stale_pdst},
     {rob_uop_1_27_stale_pdst},
     {rob_uop_1_26_stale_pdst},
     {rob_uop_1_25_stale_pdst},
     {rob_uop_1_24_stale_pdst},
     {rob_uop_1_23_stale_pdst},
     {rob_uop_1_22_stale_pdst},
     {rob_uop_1_21_stale_pdst},
     {rob_uop_1_20_stale_pdst},
     {rob_uop_1_19_stale_pdst},
     {rob_uop_1_18_stale_pdst},
     {rob_uop_1_17_stale_pdst},
     {rob_uop_1_16_stale_pdst},
     {rob_uop_1_15_stale_pdst},
     {rob_uop_1_14_stale_pdst},
     {rob_uop_1_13_stale_pdst},
     {rob_uop_1_12_stale_pdst},
     {rob_uop_1_11_stale_pdst},
     {rob_uop_1_10_stale_pdst},
     {rob_uop_1_9_stale_pdst},
     {rob_uop_1_8_stale_pdst},
     {rob_uop_1_7_stale_pdst},
     {rob_uop_1_6_stale_pdst},
     {rob_uop_1_5_stale_pdst},
     {rob_uop_1_4_stale_pdst},
     {rob_uop_1_3_stale_pdst},
     {rob_uop_1_2_stale_pdst},
     {rob_uop_1_1_stale_pdst},
     {rob_uop_1_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_50 =
    {{rob_uop_1_31_is_fencei},
     {rob_uop_1_30_is_fencei},
     {rob_uop_1_29_is_fencei},
     {rob_uop_1_28_is_fencei},
     {rob_uop_1_27_is_fencei},
     {rob_uop_1_26_is_fencei},
     {rob_uop_1_25_is_fencei},
     {rob_uop_1_24_is_fencei},
     {rob_uop_1_23_is_fencei},
     {rob_uop_1_22_is_fencei},
     {rob_uop_1_21_is_fencei},
     {rob_uop_1_20_is_fencei},
     {rob_uop_1_19_is_fencei},
     {rob_uop_1_18_is_fencei},
     {rob_uop_1_17_is_fencei},
     {rob_uop_1_16_is_fencei},
     {rob_uop_1_15_is_fencei},
     {rob_uop_1_14_is_fencei},
     {rob_uop_1_13_is_fencei},
     {rob_uop_1_12_is_fencei},
     {rob_uop_1_11_is_fencei},
     {rob_uop_1_10_is_fencei},
     {rob_uop_1_9_is_fencei},
     {rob_uop_1_8_is_fencei},
     {rob_uop_1_7_is_fencei},
     {rob_uop_1_6_is_fencei},
     {rob_uop_1_5_is_fencei},
     {rob_uop_1_4_is_fencei},
     {rob_uop_1_3_is_fencei},
     {rob_uop_1_2_is_fencei},
     {rob_uop_1_1_is_fencei},
     {rob_uop_1_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_51 =
    {{rob_uop_1_31_uses_ldq},
     {rob_uop_1_30_uses_ldq},
     {rob_uop_1_29_uses_ldq},
     {rob_uop_1_28_uses_ldq},
     {rob_uop_1_27_uses_ldq},
     {rob_uop_1_26_uses_ldq},
     {rob_uop_1_25_uses_ldq},
     {rob_uop_1_24_uses_ldq},
     {rob_uop_1_23_uses_ldq},
     {rob_uop_1_22_uses_ldq},
     {rob_uop_1_21_uses_ldq},
     {rob_uop_1_20_uses_ldq},
     {rob_uop_1_19_uses_ldq},
     {rob_uop_1_18_uses_ldq},
     {rob_uop_1_17_uses_ldq},
     {rob_uop_1_16_uses_ldq},
     {rob_uop_1_15_uses_ldq},
     {rob_uop_1_14_uses_ldq},
     {rob_uop_1_13_uses_ldq},
     {rob_uop_1_12_uses_ldq},
     {rob_uop_1_11_uses_ldq},
     {rob_uop_1_10_uses_ldq},
     {rob_uop_1_9_uses_ldq},
     {rob_uop_1_8_uses_ldq},
     {rob_uop_1_7_uses_ldq},
     {rob_uop_1_6_uses_ldq},
     {rob_uop_1_5_uses_ldq},
     {rob_uop_1_4_uses_ldq},
     {rob_uop_1_3_uses_ldq},
     {rob_uop_1_2_uses_ldq},
     {rob_uop_1_1_uses_ldq},
     {rob_uop_1_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_52 =
    {{rob_uop_1_31_uses_stq},
     {rob_uop_1_30_uses_stq},
     {rob_uop_1_29_uses_stq},
     {rob_uop_1_28_uses_stq},
     {rob_uop_1_27_uses_stq},
     {rob_uop_1_26_uses_stq},
     {rob_uop_1_25_uses_stq},
     {rob_uop_1_24_uses_stq},
     {rob_uop_1_23_uses_stq},
     {rob_uop_1_22_uses_stq},
     {rob_uop_1_21_uses_stq},
     {rob_uop_1_20_uses_stq},
     {rob_uop_1_19_uses_stq},
     {rob_uop_1_18_uses_stq},
     {rob_uop_1_17_uses_stq},
     {rob_uop_1_16_uses_stq},
     {rob_uop_1_15_uses_stq},
     {rob_uop_1_14_uses_stq},
     {rob_uop_1_13_uses_stq},
     {rob_uop_1_12_uses_stq},
     {rob_uop_1_11_uses_stq},
     {rob_uop_1_10_uses_stq},
     {rob_uop_1_9_uses_stq},
     {rob_uop_1_8_uses_stq},
     {rob_uop_1_7_uses_stq},
     {rob_uop_1_6_uses_stq},
     {rob_uop_1_5_uses_stq},
     {rob_uop_1_4_uses_stq},
     {rob_uop_1_3_uses_stq},
     {rob_uop_1_2_uses_stq},
     {rob_uop_1_1_uses_stq},
     {rob_uop_1_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_53 =
    {{rob_uop_1_31_is_sys_pc2epc},
     {rob_uop_1_30_is_sys_pc2epc},
     {rob_uop_1_29_is_sys_pc2epc},
     {rob_uop_1_28_is_sys_pc2epc},
     {rob_uop_1_27_is_sys_pc2epc},
     {rob_uop_1_26_is_sys_pc2epc},
     {rob_uop_1_25_is_sys_pc2epc},
     {rob_uop_1_24_is_sys_pc2epc},
     {rob_uop_1_23_is_sys_pc2epc},
     {rob_uop_1_22_is_sys_pc2epc},
     {rob_uop_1_21_is_sys_pc2epc},
     {rob_uop_1_20_is_sys_pc2epc},
     {rob_uop_1_19_is_sys_pc2epc},
     {rob_uop_1_18_is_sys_pc2epc},
     {rob_uop_1_17_is_sys_pc2epc},
     {rob_uop_1_16_is_sys_pc2epc},
     {rob_uop_1_15_is_sys_pc2epc},
     {rob_uop_1_14_is_sys_pc2epc},
     {rob_uop_1_13_is_sys_pc2epc},
     {rob_uop_1_12_is_sys_pc2epc},
     {rob_uop_1_11_is_sys_pc2epc},
     {rob_uop_1_10_is_sys_pc2epc},
     {rob_uop_1_9_is_sys_pc2epc},
     {rob_uop_1_8_is_sys_pc2epc},
     {rob_uop_1_7_is_sys_pc2epc},
     {rob_uop_1_6_is_sys_pc2epc},
     {rob_uop_1_5_is_sys_pc2epc},
     {rob_uop_1_4_is_sys_pc2epc},
     {rob_uop_1_3_is_sys_pc2epc},
     {rob_uop_1_2_is_sys_pc2epc},
     {rob_uop_1_1_is_sys_pc2epc},
     {rob_uop_1_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_54 =
    {{rob_uop_1_31_flush_on_commit},
     {rob_uop_1_30_flush_on_commit},
     {rob_uop_1_29_flush_on_commit},
     {rob_uop_1_28_flush_on_commit},
     {rob_uop_1_27_flush_on_commit},
     {rob_uop_1_26_flush_on_commit},
     {rob_uop_1_25_flush_on_commit},
     {rob_uop_1_24_flush_on_commit},
     {rob_uop_1_23_flush_on_commit},
     {rob_uop_1_22_flush_on_commit},
     {rob_uop_1_21_flush_on_commit},
     {rob_uop_1_20_flush_on_commit},
     {rob_uop_1_19_flush_on_commit},
     {rob_uop_1_18_flush_on_commit},
     {rob_uop_1_17_flush_on_commit},
     {rob_uop_1_16_flush_on_commit},
     {rob_uop_1_15_flush_on_commit},
     {rob_uop_1_14_flush_on_commit},
     {rob_uop_1_13_flush_on_commit},
     {rob_uop_1_12_flush_on_commit},
     {rob_uop_1_11_flush_on_commit},
     {rob_uop_1_10_flush_on_commit},
     {rob_uop_1_9_flush_on_commit},
     {rob_uop_1_8_flush_on_commit},
     {rob_uop_1_7_flush_on_commit},
     {rob_uop_1_6_flush_on_commit},
     {rob_uop_1_5_flush_on_commit},
     {rob_uop_1_4_flush_on_commit},
     {rob_uop_1_3_flush_on_commit},
     {rob_uop_1_2_flush_on_commit},
     {rob_uop_1_1_flush_on_commit},
     {rob_uop_1_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_55 =
    {{rob_uop_1_31_ldst},
     {rob_uop_1_30_ldst},
     {rob_uop_1_29_ldst},
     {rob_uop_1_28_ldst},
     {rob_uop_1_27_ldst},
     {rob_uop_1_26_ldst},
     {rob_uop_1_25_ldst},
     {rob_uop_1_24_ldst},
     {rob_uop_1_23_ldst},
     {rob_uop_1_22_ldst},
     {rob_uop_1_21_ldst},
     {rob_uop_1_20_ldst},
     {rob_uop_1_19_ldst},
     {rob_uop_1_18_ldst},
     {rob_uop_1_17_ldst},
     {rob_uop_1_16_ldst},
     {rob_uop_1_15_ldst},
     {rob_uop_1_14_ldst},
     {rob_uop_1_13_ldst},
     {rob_uop_1_12_ldst},
     {rob_uop_1_11_ldst},
     {rob_uop_1_10_ldst},
     {rob_uop_1_9_ldst},
     {rob_uop_1_8_ldst},
     {rob_uop_1_7_ldst},
     {rob_uop_1_6_ldst},
     {rob_uop_1_5_ldst},
     {rob_uop_1_4_ldst},
     {rob_uop_1_3_ldst},
     {rob_uop_1_2_ldst},
     {rob_uop_1_1_ldst},
     {rob_uop_1_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_56 =
    {{rob_uop_1_31_ldst_val},
     {rob_uop_1_30_ldst_val},
     {rob_uop_1_29_ldst_val},
     {rob_uop_1_28_ldst_val},
     {rob_uop_1_27_ldst_val},
     {rob_uop_1_26_ldst_val},
     {rob_uop_1_25_ldst_val},
     {rob_uop_1_24_ldst_val},
     {rob_uop_1_23_ldst_val},
     {rob_uop_1_22_ldst_val},
     {rob_uop_1_21_ldst_val},
     {rob_uop_1_20_ldst_val},
     {rob_uop_1_19_ldst_val},
     {rob_uop_1_18_ldst_val},
     {rob_uop_1_17_ldst_val},
     {rob_uop_1_16_ldst_val},
     {rob_uop_1_15_ldst_val},
     {rob_uop_1_14_ldst_val},
     {rob_uop_1_13_ldst_val},
     {rob_uop_1_12_ldst_val},
     {rob_uop_1_11_ldst_val},
     {rob_uop_1_10_ldst_val},
     {rob_uop_1_9_ldst_val},
     {rob_uop_1_8_ldst_val},
     {rob_uop_1_7_ldst_val},
     {rob_uop_1_6_ldst_val},
     {rob_uop_1_5_ldst_val},
     {rob_uop_1_4_ldst_val},
     {rob_uop_1_3_ldst_val},
     {rob_uop_1_2_ldst_val},
     {rob_uop_1_1_ldst_val},
     {rob_uop_1_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_57 =
    {{rob_uop_1_31_dst_rtype},
     {rob_uop_1_30_dst_rtype},
     {rob_uop_1_29_dst_rtype},
     {rob_uop_1_28_dst_rtype},
     {rob_uop_1_27_dst_rtype},
     {rob_uop_1_26_dst_rtype},
     {rob_uop_1_25_dst_rtype},
     {rob_uop_1_24_dst_rtype},
     {rob_uop_1_23_dst_rtype},
     {rob_uop_1_22_dst_rtype},
     {rob_uop_1_21_dst_rtype},
     {rob_uop_1_20_dst_rtype},
     {rob_uop_1_19_dst_rtype},
     {rob_uop_1_18_dst_rtype},
     {rob_uop_1_17_dst_rtype},
     {rob_uop_1_16_dst_rtype},
     {rob_uop_1_15_dst_rtype},
     {rob_uop_1_14_dst_rtype},
     {rob_uop_1_13_dst_rtype},
     {rob_uop_1_12_dst_rtype},
     {rob_uop_1_11_dst_rtype},
     {rob_uop_1_10_dst_rtype},
     {rob_uop_1_9_dst_rtype},
     {rob_uop_1_8_dst_rtype},
     {rob_uop_1_7_dst_rtype},
     {rob_uop_1_6_dst_rtype},
     {rob_uop_1_5_dst_rtype},
     {rob_uop_1_4_dst_rtype},
     {rob_uop_1_3_dst_rtype},
     {rob_uop_1_2_dst_rtype},
     {rob_uop_1_1_dst_rtype},
     {rob_uop_1_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_58 =
    {{rob_uop_1_31_fp_val},
     {rob_uop_1_30_fp_val},
     {rob_uop_1_29_fp_val},
     {rob_uop_1_28_fp_val},
     {rob_uop_1_27_fp_val},
     {rob_uop_1_26_fp_val},
     {rob_uop_1_25_fp_val},
     {rob_uop_1_24_fp_val},
     {rob_uop_1_23_fp_val},
     {rob_uop_1_22_fp_val},
     {rob_uop_1_21_fp_val},
     {rob_uop_1_20_fp_val},
     {rob_uop_1_19_fp_val},
     {rob_uop_1_18_fp_val},
     {rob_uop_1_17_fp_val},
     {rob_uop_1_16_fp_val},
     {rob_uop_1_15_fp_val},
     {rob_uop_1_14_fp_val},
     {rob_uop_1_13_fp_val},
     {rob_uop_1_12_fp_val},
     {rob_uop_1_11_fp_val},
     {rob_uop_1_10_fp_val},
     {rob_uop_1_9_fp_val},
     {rob_uop_1_8_fp_val},
     {rob_uop_1_7_fp_val},
     {rob_uop_1_6_fp_val},
     {rob_uop_1_5_fp_val},
     {rob_uop_1_4_fp_val},
     {rob_uop_1_3_fp_val},
     {rob_uop_1_2_fp_val},
     {rob_uop_1_1_fp_val},
     {rob_uop_1_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row_1 = _io_commit_rollback_T_2 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_1_output = rbk_row_1 & _GEN_29[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              rob_val_2_0;	// rob.scala:307:32
  reg              rob_val_2_1;	// rob.scala:307:32
  reg              rob_val_2_2;	// rob.scala:307:32
  reg              rob_val_2_3;	// rob.scala:307:32
  reg              rob_val_2_4;	// rob.scala:307:32
  reg              rob_val_2_5;	// rob.scala:307:32
  reg              rob_val_2_6;	// rob.scala:307:32
  reg              rob_val_2_7;	// rob.scala:307:32
  reg              rob_val_2_8;	// rob.scala:307:32
  reg              rob_val_2_9;	// rob.scala:307:32
  reg              rob_val_2_10;	// rob.scala:307:32
  reg              rob_val_2_11;	// rob.scala:307:32
  reg              rob_val_2_12;	// rob.scala:307:32
  reg              rob_val_2_13;	// rob.scala:307:32
  reg              rob_val_2_14;	// rob.scala:307:32
  reg              rob_val_2_15;	// rob.scala:307:32
  reg              rob_val_2_16;	// rob.scala:307:32
  reg              rob_val_2_17;	// rob.scala:307:32
  reg              rob_val_2_18;	// rob.scala:307:32
  reg              rob_val_2_19;	// rob.scala:307:32
  reg              rob_val_2_20;	// rob.scala:307:32
  reg              rob_val_2_21;	// rob.scala:307:32
  reg              rob_val_2_22;	// rob.scala:307:32
  reg              rob_val_2_23;	// rob.scala:307:32
  reg              rob_val_2_24;	// rob.scala:307:32
  reg              rob_val_2_25;	// rob.scala:307:32
  reg              rob_val_2_26;	// rob.scala:307:32
  reg              rob_val_2_27;	// rob.scala:307:32
  reg              rob_val_2_28;	// rob.scala:307:32
  reg              rob_val_2_29;	// rob.scala:307:32
  reg              rob_val_2_30;	// rob.scala:307:32
  reg              rob_val_2_31;	// rob.scala:307:32
  reg              rob_bsy_2_0;	// rob.scala:308:28
  reg              rob_bsy_2_1;	// rob.scala:308:28
  reg              rob_bsy_2_2;	// rob.scala:308:28
  reg              rob_bsy_2_3;	// rob.scala:308:28
  reg              rob_bsy_2_4;	// rob.scala:308:28
  reg              rob_bsy_2_5;	// rob.scala:308:28
  reg              rob_bsy_2_6;	// rob.scala:308:28
  reg              rob_bsy_2_7;	// rob.scala:308:28
  reg              rob_bsy_2_8;	// rob.scala:308:28
  reg              rob_bsy_2_9;	// rob.scala:308:28
  reg              rob_bsy_2_10;	// rob.scala:308:28
  reg              rob_bsy_2_11;	// rob.scala:308:28
  reg              rob_bsy_2_12;	// rob.scala:308:28
  reg              rob_bsy_2_13;	// rob.scala:308:28
  reg              rob_bsy_2_14;	// rob.scala:308:28
  reg              rob_bsy_2_15;	// rob.scala:308:28
  reg              rob_bsy_2_16;	// rob.scala:308:28
  reg              rob_bsy_2_17;	// rob.scala:308:28
  reg              rob_bsy_2_18;	// rob.scala:308:28
  reg              rob_bsy_2_19;	// rob.scala:308:28
  reg              rob_bsy_2_20;	// rob.scala:308:28
  reg              rob_bsy_2_21;	// rob.scala:308:28
  reg              rob_bsy_2_22;	// rob.scala:308:28
  reg              rob_bsy_2_23;	// rob.scala:308:28
  reg              rob_bsy_2_24;	// rob.scala:308:28
  reg              rob_bsy_2_25;	// rob.scala:308:28
  reg              rob_bsy_2_26;	// rob.scala:308:28
  reg              rob_bsy_2_27;	// rob.scala:308:28
  reg              rob_bsy_2_28;	// rob.scala:308:28
  reg              rob_bsy_2_29;	// rob.scala:308:28
  reg              rob_bsy_2_30;	// rob.scala:308:28
  reg              rob_bsy_2_31;	// rob.scala:308:28
  reg              rob_unsafe_2_0;	// rob.scala:309:28
  reg              rob_unsafe_2_1;	// rob.scala:309:28
  reg              rob_unsafe_2_2;	// rob.scala:309:28
  reg              rob_unsafe_2_3;	// rob.scala:309:28
  reg              rob_unsafe_2_4;	// rob.scala:309:28
  reg              rob_unsafe_2_5;	// rob.scala:309:28
  reg              rob_unsafe_2_6;	// rob.scala:309:28
  reg              rob_unsafe_2_7;	// rob.scala:309:28
  reg              rob_unsafe_2_8;	// rob.scala:309:28
  reg              rob_unsafe_2_9;	// rob.scala:309:28
  reg              rob_unsafe_2_10;	// rob.scala:309:28
  reg              rob_unsafe_2_11;	// rob.scala:309:28
  reg              rob_unsafe_2_12;	// rob.scala:309:28
  reg              rob_unsafe_2_13;	// rob.scala:309:28
  reg              rob_unsafe_2_14;	// rob.scala:309:28
  reg              rob_unsafe_2_15;	// rob.scala:309:28
  reg              rob_unsafe_2_16;	// rob.scala:309:28
  reg              rob_unsafe_2_17;	// rob.scala:309:28
  reg              rob_unsafe_2_18;	// rob.scala:309:28
  reg              rob_unsafe_2_19;	// rob.scala:309:28
  reg              rob_unsafe_2_20;	// rob.scala:309:28
  reg              rob_unsafe_2_21;	// rob.scala:309:28
  reg              rob_unsafe_2_22;	// rob.scala:309:28
  reg              rob_unsafe_2_23;	// rob.scala:309:28
  reg              rob_unsafe_2_24;	// rob.scala:309:28
  reg              rob_unsafe_2_25;	// rob.scala:309:28
  reg              rob_unsafe_2_26;	// rob.scala:309:28
  reg              rob_unsafe_2_27;	// rob.scala:309:28
  reg              rob_unsafe_2_28;	// rob.scala:309:28
  reg              rob_unsafe_2_29;	// rob.scala:309:28
  reg              rob_unsafe_2_30;	// rob.scala:309:28
  reg              rob_unsafe_2_31;	// rob.scala:309:28
  reg  [6:0]       rob_uop_2_0_uopc;	// rob.scala:310:28
  reg              rob_uop_2_0_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_0_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_0_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_0_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_0_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_0_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_0_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_0_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_0_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_0_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_0_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_0_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_0_ldst;	// rob.scala:310:28
  reg              rob_uop_2_0_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_0_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_0_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_1_uopc;	// rob.scala:310:28
  reg              rob_uop_2_1_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_1_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_1_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_1_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_1_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_1_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_1_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_1_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_1_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_1_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_1_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_1_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_1_ldst;	// rob.scala:310:28
  reg              rob_uop_2_1_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_1_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_1_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_2_uopc;	// rob.scala:310:28
  reg              rob_uop_2_2_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_2_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_2_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_2_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_2_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_2_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_2_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_2_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_2_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_2_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_2_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_2_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_2_ldst;	// rob.scala:310:28
  reg              rob_uop_2_2_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_2_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_2_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_3_uopc;	// rob.scala:310:28
  reg              rob_uop_2_3_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_3_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_3_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_3_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_3_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_3_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_3_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_3_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_3_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_3_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_3_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_3_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_3_ldst;	// rob.scala:310:28
  reg              rob_uop_2_3_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_3_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_3_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_4_uopc;	// rob.scala:310:28
  reg              rob_uop_2_4_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_4_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_4_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_4_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_4_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_4_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_4_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_4_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_4_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_4_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_4_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_4_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_4_ldst;	// rob.scala:310:28
  reg              rob_uop_2_4_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_4_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_4_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_5_uopc;	// rob.scala:310:28
  reg              rob_uop_2_5_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_5_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_5_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_5_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_5_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_5_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_5_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_5_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_5_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_5_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_5_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_5_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_5_ldst;	// rob.scala:310:28
  reg              rob_uop_2_5_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_5_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_5_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_6_uopc;	// rob.scala:310:28
  reg              rob_uop_2_6_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_6_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_6_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_6_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_6_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_6_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_6_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_6_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_6_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_6_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_6_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_6_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_6_ldst;	// rob.scala:310:28
  reg              rob_uop_2_6_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_6_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_6_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_7_uopc;	// rob.scala:310:28
  reg              rob_uop_2_7_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_7_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_7_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_7_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_7_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_7_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_7_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_7_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_7_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_7_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_7_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_7_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_7_ldst;	// rob.scala:310:28
  reg              rob_uop_2_7_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_7_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_7_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_8_uopc;	// rob.scala:310:28
  reg              rob_uop_2_8_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_8_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_8_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_8_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_8_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_8_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_8_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_8_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_8_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_8_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_8_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_8_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_8_ldst;	// rob.scala:310:28
  reg              rob_uop_2_8_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_8_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_8_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_9_uopc;	// rob.scala:310:28
  reg              rob_uop_2_9_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_9_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_9_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_9_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_9_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_9_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_9_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_9_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_9_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_9_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_9_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_9_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_9_ldst;	// rob.scala:310:28
  reg              rob_uop_2_9_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_9_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_9_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_10_uopc;	// rob.scala:310:28
  reg              rob_uop_2_10_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_10_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_10_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_10_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_10_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_10_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_10_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_10_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_10_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_10_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_10_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_10_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_10_ldst;	// rob.scala:310:28
  reg              rob_uop_2_10_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_10_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_10_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_11_uopc;	// rob.scala:310:28
  reg              rob_uop_2_11_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_11_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_11_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_11_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_11_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_11_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_11_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_11_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_11_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_11_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_11_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_11_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_11_ldst;	// rob.scala:310:28
  reg              rob_uop_2_11_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_11_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_11_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_12_uopc;	// rob.scala:310:28
  reg              rob_uop_2_12_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_12_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_12_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_12_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_12_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_12_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_12_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_12_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_12_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_12_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_12_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_12_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_12_ldst;	// rob.scala:310:28
  reg              rob_uop_2_12_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_12_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_12_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_13_uopc;	// rob.scala:310:28
  reg              rob_uop_2_13_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_13_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_13_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_13_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_13_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_13_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_13_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_13_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_13_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_13_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_13_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_13_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_13_ldst;	// rob.scala:310:28
  reg              rob_uop_2_13_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_13_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_13_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_14_uopc;	// rob.scala:310:28
  reg              rob_uop_2_14_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_14_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_14_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_14_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_14_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_14_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_14_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_14_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_14_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_14_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_14_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_14_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_14_ldst;	// rob.scala:310:28
  reg              rob_uop_2_14_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_14_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_14_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_15_uopc;	// rob.scala:310:28
  reg              rob_uop_2_15_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_15_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_15_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_15_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_15_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_15_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_15_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_15_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_15_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_15_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_15_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_15_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_15_ldst;	// rob.scala:310:28
  reg              rob_uop_2_15_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_15_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_15_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_16_uopc;	// rob.scala:310:28
  reg              rob_uop_2_16_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_16_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_16_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_16_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_16_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_16_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_16_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_16_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_16_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_16_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_16_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_16_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_16_ldst;	// rob.scala:310:28
  reg              rob_uop_2_16_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_16_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_16_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_17_uopc;	// rob.scala:310:28
  reg              rob_uop_2_17_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_17_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_17_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_17_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_17_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_17_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_17_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_17_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_17_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_17_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_17_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_17_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_17_ldst;	// rob.scala:310:28
  reg              rob_uop_2_17_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_17_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_17_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_18_uopc;	// rob.scala:310:28
  reg              rob_uop_2_18_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_18_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_18_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_18_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_18_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_18_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_18_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_18_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_18_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_18_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_18_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_18_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_18_ldst;	// rob.scala:310:28
  reg              rob_uop_2_18_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_18_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_18_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_19_uopc;	// rob.scala:310:28
  reg              rob_uop_2_19_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_19_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_19_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_19_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_19_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_19_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_19_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_19_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_19_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_19_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_19_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_19_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_19_ldst;	// rob.scala:310:28
  reg              rob_uop_2_19_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_19_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_19_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_20_uopc;	// rob.scala:310:28
  reg              rob_uop_2_20_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_20_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_20_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_20_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_20_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_20_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_20_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_20_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_20_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_20_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_20_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_20_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_20_ldst;	// rob.scala:310:28
  reg              rob_uop_2_20_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_20_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_20_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_21_uopc;	// rob.scala:310:28
  reg              rob_uop_2_21_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_21_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_21_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_21_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_21_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_21_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_21_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_21_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_21_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_21_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_21_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_21_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_21_ldst;	// rob.scala:310:28
  reg              rob_uop_2_21_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_21_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_21_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_22_uopc;	// rob.scala:310:28
  reg              rob_uop_2_22_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_22_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_22_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_22_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_22_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_22_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_22_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_22_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_22_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_22_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_22_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_22_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_22_ldst;	// rob.scala:310:28
  reg              rob_uop_2_22_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_22_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_22_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_23_uopc;	// rob.scala:310:28
  reg              rob_uop_2_23_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_23_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_23_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_23_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_23_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_23_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_23_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_23_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_23_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_23_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_23_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_23_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_23_ldst;	// rob.scala:310:28
  reg              rob_uop_2_23_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_23_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_23_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_24_uopc;	// rob.scala:310:28
  reg              rob_uop_2_24_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_24_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_24_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_24_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_24_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_24_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_24_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_24_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_24_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_24_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_24_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_24_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_24_ldst;	// rob.scala:310:28
  reg              rob_uop_2_24_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_24_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_24_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_25_uopc;	// rob.scala:310:28
  reg              rob_uop_2_25_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_25_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_25_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_25_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_25_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_25_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_25_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_25_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_25_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_25_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_25_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_25_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_25_ldst;	// rob.scala:310:28
  reg              rob_uop_2_25_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_25_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_25_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_26_uopc;	// rob.scala:310:28
  reg              rob_uop_2_26_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_26_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_26_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_26_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_26_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_26_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_26_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_26_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_26_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_26_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_26_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_26_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_26_ldst;	// rob.scala:310:28
  reg              rob_uop_2_26_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_26_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_26_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_27_uopc;	// rob.scala:310:28
  reg              rob_uop_2_27_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_27_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_27_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_27_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_27_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_27_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_27_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_27_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_27_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_27_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_27_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_27_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_27_ldst;	// rob.scala:310:28
  reg              rob_uop_2_27_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_27_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_27_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_28_uopc;	// rob.scala:310:28
  reg              rob_uop_2_28_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_28_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_28_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_28_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_28_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_28_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_28_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_28_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_28_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_28_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_28_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_28_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_28_ldst;	// rob.scala:310:28
  reg              rob_uop_2_28_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_28_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_28_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_29_uopc;	// rob.scala:310:28
  reg              rob_uop_2_29_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_29_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_29_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_29_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_29_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_29_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_29_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_29_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_29_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_29_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_29_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_29_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_29_ldst;	// rob.scala:310:28
  reg              rob_uop_2_29_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_29_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_29_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_30_uopc;	// rob.scala:310:28
  reg              rob_uop_2_30_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_30_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_30_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_30_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_30_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_30_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_30_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_30_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_30_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_30_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_30_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_30_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_30_ldst;	// rob.scala:310:28
  reg              rob_uop_2_30_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_30_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_30_fp_val;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_31_uopc;	// rob.scala:310:28
  reg              rob_uop_2_31_is_rvc;	// rob.scala:310:28
  reg  [15:0]      rob_uop_2_31_br_mask;	// rob.scala:310:28
  reg  [4:0]       rob_uop_2_31_ftq_idx;	// rob.scala:310:28
  reg              rob_uop_2_31_edge_inst;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_31_pc_lob;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_31_pdst;	// rob.scala:310:28
  reg  [6:0]       rob_uop_2_31_stale_pdst;	// rob.scala:310:28
  reg              rob_uop_2_31_is_fencei;	// rob.scala:310:28
  reg              rob_uop_2_31_uses_ldq;	// rob.scala:310:28
  reg              rob_uop_2_31_uses_stq;	// rob.scala:310:28
  reg              rob_uop_2_31_is_sys_pc2epc;	// rob.scala:310:28
  reg              rob_uop_2_31_flush_on_commit;	// rob.scala:310:28
  reg  [5:0]       rob_uop_2_31_ldst;	// rob.scala:310:28
  reg              rob_uop_2_31_ldst_val;	// rob.scala:310:28
  reg  [1:0]       rob_uop_2_31_dst_rtype;	// rob.scala:310:28
  reg              rob_uop_2_31_fp_val;	// rob.scala:310:28
  reg              rob_exception_2_0;	// rob.scala:311:28
  reg              rob_exception_2_1;	// rob.scala:311:28
  reg              rob_exception_2_2;	// rob.scala:311:28
  reg              rob_exception_2_3;	// rob.scala:311:28
  reg              rob_exception_2_4;	// rob.scala:311:28
  reg              rob_exception_2_5;	// rob.scala:311:28
  reg              rob_exception_2_6;	// rob.scala:311:28
  reg              rob_exception_2_7;	// rob.scala:311:28
  reg              rob_exception_2_8;	// rob.scala:311:28
  reg              rob_exception_2_9;	// rob.scala:311:28
  reg              rob_exception_2_10;	// rob.scala:311:28
  reg              rob_exception_2_11;	// rob.scala:311:28
  reg              rob_exception_2_12;	// rob.scala:311:28
  reg              rob_exception_2_13;	// rob.scala:311:28
  reg              rob_exception_2_14;	// rob.scala:311:28
  reg              rob_exception_2_15;	// rob.scala:311:28
  reg              rob_exception_2_16;	// rob.scala:311:28
  reg              rob_exception_2_17;	// rob.scala:311:28
  reg              rob_exception_2_18;	// rob.scala:311:28
  reg              rob_exception_2_19;	// rob.scala:311:28
  reg              rob_exception_2_20;	// rob.scala:311:28
  reg              rob_exception_2_21;	// rob.scala:311:28
  reg              rob_exception_2_22;	// rob.scala:311:28
  reg              rob_exception_2_23;	// rob.scala:311:28
  reg              rob_exception_2_24;	// rob.scala:311:28
  reg              rob_exception_2_25;	// rob.scala:311:28
  reg              rob_exception_2_26;	// rob.scala:311:28
  reg              rob_exception_2_27;	// rob.scala:311:28
  reg              rob_exception_2_28;	// rob.scala:311:28
  reg              rob_exception_2_29;	// rob.scala:311:28
  reg              rob_exception_2_30;	// rob.scala:311:28
  reg              rob_exception_2_31;	// rob.scala:311:28
  reg              rob_predicated_2_0;	// rob.scala:312:29
  reg              rob_predicated_2_1;	// rob.scala:312:29
  reg              rob_predicated_2_2;	// rob.scala:312:29
  reg              rob_predicated_2_3;	// rob.scala:312:29
  reg              rob_predicated_2_4;	// rob.scala:312:29
  reg              rob_predicated_2_5;	// rob.scala:312:29
  reg              rob_predicated_2_6;	// rob.scala:312:29
  reg              rob_predicated_2_7;	// rob.scala:312:29
  reg              rob_predicated_2_8;	// rob.scala:312:29
  reg              rob_predicated_2_9;	// rob.scala:312:29
  reg              rob_predicated_2_10;	// rob.scala:312:29
  reg              rob_predicated_2_11;	// rob.scala:312:29
  reg              rob_predicated_2_12;	// rob.scala:312:29
  reg              rob_predicated_2_13;	// rob.scala:312:29
  reg              rob_predicated_2_14;	// rob.scala:312:29
  reg              rob_predicated_2_15;	// rob.scala:312:29
  reg              rob_predicated_2_16;	// rob.scala:312:29
  reg              rob_predicated_2_17;	// rob.scala:312:29
  reg              rob_predicated_2_18;	// rob.scala:312:29
  reg              rob_predicated_2_19;	// rob.scala:312:29
  reg              rob_predicated_2_20;	// rob.scala:312:29
  reg              rob_predicated_2_21;	// rob.scala:312:29
  reg              rob_predicated_2_22;	// rob.scala:312:29
  reg              rob_predicated_2_23;	// rob.scala:312:29
  reg              rob_predicated_2_24;	// rob.scala:312:29
  reg              rob_predicated_2_25;	// rob.scala:312:29
  reg              rob_predicated_2_26;	// rob.scala:312:29
  reg              rob_predicated_2_27;	// rob.scala:312:29
  reg              rob_predicated_2_28;	// rob.scala:312:29
  reg              rob_predicated_2_29;	// rob.scala:312:29
  reg              rob_predicated_2_30;	// rob.scala:312:29
  reg              rob_predicated_2_31;	// rob.scala:312:29
  wire [31:0]      _GEN_59 =
    {{rob_val_2_31},
     {rob_val_2_30},
     {rob_val_2_29},
     {rob_val_2_28},
     {rob_val_2_27},
     {rob_val_2_26},
     {rob_val_2_25},
     {rob_val_2_24},
     {rob_val_2_23},
     {rob_val_2_22},
     {rob_val_2_21},
     {rob_val_2_20},
     {rob_val_2_19},
     {rob_val_2_18},
     {rob_val_2_17},
     {rob_val_2_16},
     {rob_val_2_15},
     {rob_val_2_14},
     {rob_val_2_13},
     {rob_val_2_12},
     {rob_val_2_11},
     {rob_val_2_10},
     {rob_val_2_9},
     {rob_val_2_8},
     {rob_val_2_7},
     {rob_val_2_6},
     {rob_val_2_5},
     {rob_val_2_4},
     {rob_val_2_3},
     {rob_val_2_2},
     {rob_val_2_1},
     {rob_val_2_0}};	// rob.scala:307:32, :324:31
  wire             rob_tail_vals_2 = _GEN_59[rob_tail];	// rob.scala:228:29, :324:31
  wire             _GEN_60 =
    io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_61 =
    io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_62 =
    io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_63 =
    io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_64 =
    io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_65 =
    io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :346:27
  wire             _GEN_66 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :361:31
  wire [31:0]      _GEN_67 =
    {{rob_bsy_2_31},
     {rob_bsy_2_30},
     {rob_bsy_2_29},
     {rob_bsy_2_28},
     {rob_bsy_2_27},
     {rob_bsy_2_26},
     {rob_bsy_2_25},
     {rob_bsy_2_24},
     {rob_bsy_2_23},
     {rob_bsy_2_22},
     {rob_bsy_2_21},
     {rob_bsy_2_20},
     {rob_bsy_2_19},
     {rob_bsy_2_18},
     {rob_bsy_2_17},
     {rob_bsy_2_16},
     {rob_bsy_2_15},
     {rob_bsy_2_14},
     {rob_bsy_2_13},
     {rob_bsy_2_12},
     {rob_bsy_2_11},
     {rob_bsy_2_10},
     {rob_bsy_2_9},
     {rob_bsy_2_8},
     {rob_bsy_2_7},
     {rob_bsy_2_6},
     {rob_bsy_2_5},
     {rob_bsy_2_4},
     {rob_bsy_2_3},
     {rob_bsy_2_2},
     {rob_bsy_2_1},
     {rob_bsy_2_0}};	// rob.scala:308:28, :366:31
  wire             _GEN_68 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :361:31
  wire             _GEN_69 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h2;	// rob.scala:236:31, :272:36, :304:53, :390:26
  wire [31:0]      _GEN_70 =
    {{rob_unsafe_2_31},
     {rob_unsafe_2_30},
     {rob_unsafe_2_29},
     {rob_unsafe_2_28},
     {rob_unsafe_2_27},
     {rob_unsafe_2_26},
     {rob_unsafe_2_25},
     {rob_unsafe_2_24},
     {rob_unsafe_2_23},
     {rob_unsafe_2_22},
     {rob_unsafe_2_21},
     {rob_unsafe_2_20},
     {rob_unsafe_2_19},
     {rob_unsafe_2_18},
     {rob_unsafe_2_17},
     {rob_unsafe_2_16},
     {rob_unsafe_2_15},
     {rob_unsafe_2_14},
     {rob_unsafe_2_13},
     {rob_unsafe_2_12},
     {rob_unsafe_2_11},
     {rob_unsafe_2_10},
     {rob_unsafe_2_9},
     {rob_unsafe_2_8},
     {rob_unsafe_2_7},
     {rob_unsafe_2_6},
     {rob_unsafe_2_5},
     {rob_unsafe_2_4},
     {rob_unsafe_2_3},
     {rob_unsafe_2_2},
     {rob_unsafe_2_1},
     {rob_unsafe_2_0}};	// rob.scala:309:28, :394:15
  wire             rob_head_vals_2 = _GEN_59[rob_head];	// rob.scala:224:29, :324:31, :398:49
  wire [31:0]      _GEN_71 =
    {{rob_exception_2_31},
     {rob_exception_2_30},
     {rob_exception_2_29},
     {rob_exception_2_28},
     {rob_exception_2_27},
     {rob_exception_2_26},
     {rob_exception_2_25},
     {rob_exception_2_24},
     {rob_exception_2_23},
     {rob_exception_2_22},
     {rob_exception_2_21},
     {rob_exception_2_20},
     {rob_exception_2_19},
     {rob_exception_2_18},
     {rob_exception_2_17},
     {rob_exception_2_16},
     {rob_exception_2_15},
     {rob_exception_2_14},
     {rob_exception_2_13},
     {rob_exception_2_12},
     {rob_exception_2_11},
     {rob_exception_2_10},
     {rob_exception_2_9},
     {rob_exception_2_8},
     {rob_exception_2_7},
     {rob_exception_2_6},
     {rob_exception_2_5},
     {rob_exception_2_4},
     {rob_exception_2_3},
     {rob_exception_2_2},
     {rob_exception_2_1},
     {rob_exception_2_0}};	// rob.scala:311:28, :398:49
  wire             can_throw_exception_2 = rob_head_vals_2 & _GEN_71[rob_head];	// rob.scala:224:29, :398:49
  wire [31:0]      _GEN_72 =
    {{rob_predicated_2_31},
     {rob_predicated_2_30},
     {rob_predicated_2_29},
     {rob_predicated_2_28},
     {rob_predicated_2_27},
     {rob_predicated_2_26},
     {rob_predicated_2_25},
     {rob_predicated_2_24},
     {rob_predicated_2_23},
     {rob_predicated_2_22},
     {rob_predicated_2_21},
     {rob_predicated_2_20},
     {rob_predicated_2_19},
     {rob_predicated_2_18},
     {rob_predicated_2_17},
     {rob_predicated_2_16},
     {rob_predicated_2_15},
     {rob_predicated_2_14},
     {rob_predicated_2_13},
     {rob_predicated_2_12},
     {rob_predicated_2_11},
     {rob_predicated_2_10},
     {rob_predicated_2_9},
     {rob_predicated_2_8},
     {rob_predicated_2_7},
     {rob_predicated_2_6},
     {rob_predicated_2_5},
     {rob_predicated_2_4},
     {rob_predicated_2_3},
     {rob_predicated_2_2},
     {rob_predicated_2_1},
     {rob_predicated_2_0}};	// rob.scala:312:29, :410:51
  wire [31:0][6:0] _GEN_73 =
    {{rob_uop_2_31_uopc},
     {rob_uop_2_30_uopc},
     {rob_uop_2_29_uopc},
     {rob_uop_2_28_uopc},
     {rob_uop_2_27_uopc},
     {rob_uop_2_26_uopc},
     {rob_uop_2_25_uopc},
     {rob_uop_2_24_uopc},
     {rob_uop_2_23_uopc},
     {rob_uop_2_22_uopc},
     {rob_uop_2_21_uopc},
     {rob_uop_2_20_uopc},
     {rob_uop_2_19_uopc},
     {rob_uop_2_18_uopc},
     {rob_uop_2_17_uopc},
     {rob_uop_2_16_uopc},
     {rob_uop_2_15_uopc},
     {rob_uop_2_14_uopc},
     {rob_uop_2_13_uopc},
     {rob_uop_2_12_uopc},
     {rob_uop_2_11_uopc},
     {rob_uop_2_10_uopc},
     {rob_uop_2_9_uopc},
     {rob_uop_2_8_uopc},
     {rob_uop_2_7_uopc},
     {rob_uop_2_6_uopc},
     {rob_uop_2_5_uopc},
     {rob_uop_2_4_uopc},
     {rob_uop_2_3_uopc},
     {rob_uop_2_2_uopc},
     {rob_uop_2_1_uopc},
     {rob_uop_2_0_uopc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_74 =
    {{rob_uop_2_31_is_rvc},
     {rob_uop_2_30_is_rvc},
     {rob_uop_2_29_is_rvc},
     {rob_uop_2_28_is_rvc},
     {rob_uop_2_27_is_rvc},
     {rob_uop_2_26_is_rvc},
     {rob_uop_2_25_is_rvc},
     {rob_uop_2_24_is_rvc},
     {rob_uop_2_23_is_rvc},
     {rob_uop_2_22_is_rvc},
     {rob_uop_2_21_is_rvc},
     {rob_uop_2_20_is_rvc},
     {rob_uop_2_19_is_rvc},
     {rob_uop_2_18_is_rvc},
     {rob_uop_2_17_is_rvc},
     {rob_uop_2_16_is_rvc},
     {rob_uop_2_15_is_rvc},
     {rob_uop_2_14_is_rvc},
     {rob_uop_2_13_is_rvc},
     {rob_uop_2_12_is_rvc},
     {rob_uop_2_11_is_rvc},
     {rob_uop_2_10_is_rvc},
     {rob_uop_2_9_is_rvc},
     {rob_uop_2_8_is_rvc},
     {rob_uop_2_7_is_rvc},
     {rob_uop_2_6_is_rvc},
     {rob_uop_2_5_is_rvc},
     {rob_uop_2_4_is_rvc},
     {rob_uop_2_3_is_rvc},
     {rob_uop_2_2_is_rvc},
     {rob_uop_2_1_is_rvc},
     {rob_uop_2_0_is_rvc}};	// rob.scala:310:28, :411:25
  wire [31:0][4:0] _GEN_75 =
    {{rob_uop_2_31_ftq_idx},
     {rob_uop_2_30_ftq_idx},
     {rob_uop_2_29_ftq_idx},
     {rob_uop_2_28_ftq_idx},
     {rob_uop_2_27_ftq_idx},
     {rob_uop_2_26_ftq_idx},
     {rob_uop_2_25_ftq_idx},
     {rob_uop_2_24_ftq_idx},
     {rob_uop_2_23_ftq_idx},
     {rob_uop_2_22_ftq_idx},
     {rob_uop_2_21_ftq_idx},
     {rob_uop_2_20_ftq_idx},
     {rob_uop_2_19_ftq_idx},
     {rob_uop_2_18_ftq_idx},
     {rob_uop_2_17_ftq_idx},
     {rob_uop_2_16_ftq_idx},
     {rob_uop_2_15_ftq_idx},
     {rob_uop_2_14_ftq_idx},
     {rob_uop_2_13_ftq_idx},
     {rob_uop_2_12_ftq_idx},
     {rob_uop_2_11_ftq_idx},
     {rob_uop_2_10_ftq_idx},
     {rob_uop_2_9_ftq_idx},
     {rob_uop_2_8_ftq_idx},
     {rob_uop_2_7_ftq_idx},
     {rob_uop_2_6_ftq_idx},
     {rob_uop_2_5_ftq_idx},
     {rob_uop_2_4_ftq_idx},
     {rob_uop_2_3_ftq_idx},
     {rob_uop_2_2_ftq_idx},
     {rob_uop_2_1_ftq_idx},
     {rob_uop_2_0_ftq_idx}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_76 =
    {{rob_uop_2_31_edge_inst},
     {rob_uop_2_30_edge_inst},
     {rob_uop_2_29_edge_inst},
     {rob_uop_2_28_edge_inst},
     {rob_uop_2_27_edge_inst},
     {rob_uop_2_26_edge_inst},
     {rob_uop_2_25_edge_inst},
     {rob_uop_2_24_edge_inst},
     {rob_uop_2_23_edge_inst},
     {rob_uop_2_22_edge_inst},
     {rob_uop_2_21_edge_inst},
     {rob_uop_2_20_edge_inst},
     {rob_uop_2_19_edge_inst},
     {rob_uop_2_18_edge_inst},
     {rob_uop_2_17_edge_inst},
     {rob_uop_2_16_edge_inst},
     {rob_uop_2_15_edge_inst},
     {rob_uop_2_14_edge_inst},
     {rob_uop_2_13_edge_inst},
     {rob_uop_2_12_edge_inst},
     {rob_uop_2_11_edge_inst},
     {rob_uop_2_10_edge_inst},
     {rob_uop_2_9_edge_inst},
     {rob_uop_2_8_edge_inst},
     {rob_uop_2_7_edge_inst},
     {rob_uop_2_6_edge_inst},
     {rob_uop_2_5_edge_inst},
     {rob_uop_2_4_edge_inst},
     {rob_uop_2_3_edge_inst},
     {rob_uop_2_2_edge_inst},
     {rob_uop_2_1_edge_inst},
     {rob_uop_2_0_edge_inst}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_77 =
    {{rob_uop_2_31_pc_lob},
     {rob_uop_2_30_pc_lob},
     {rob_uop_2_29_pc_lob},
     {rob_uop_2_28_pc_lob},
     {rob_uop_2_27_pc_lob},
     {rob_uop_2_26_pc_lob},
     {rob_uop_2_25_pc_lob},
     {rob_uop_2_24_pc_lob},
     {rob_uop_2_23_pc_lob},
     {rob_uop_2_22_pc_lob},
     {rob_uop_2_21_pc_lob},
     {rob_uop_2_20_pc_lob},
     {rob_uop_2_19_pc_lob},
     {rob_uop_2_18_pc_lob},
     {rob_uop_2_17_pc_lob},
     {rob_uop_2_16_pc_lob},
     {rob_uop_2_15_pc_lob},
     {rob_uop_2_14_pc_lob},
     {rob_uop_2_13_pc_lob},
     {rob_uop_2_12_pc_lob},
     {rob_uop_2_11_pc_lob},
     {rob_uop_2_10_pc_lob},
     {rob_uop_2_9_pc_lob},
     {rob_uop_2_8_pc_lob},
     {rob_uop_2_7_pc_lob},
     {rob_uop_2_6_pc_lob},
     {rob_uop_2_5_pc_lob},
     {rob_uop_2_4_pc_lob},
     {rob_uop_2_3_pc_lob},
     {rob_uop_2_2_pc_lob},
     {rob_uop_2_1_pc_lob},
     {rob_uop_2_0_pc_lob}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_78 =
    {{rob_uop_2_31_pdst},
     {rob_uop_2_30_pdst},
     {rob_uop_2_29_pdst},
     {rob_uop_2_28_pdst},
     {rob_uop_2_27_pdst},
     {rob_uop_2_26_pdst},
     {rob_uop_2_25_pdst},
     {rob_uop_2_24_pdst},
     {rob_uop_2_23_pdst},
     {rob_uop_2_22_pdst},
     {rob_uop_2_21_pdst},
     {rob_uop_2_20_pdst},
     {rob_uop_2_19_pdst},
     {rob_uop_2_18_pdst},
     {rob_uop_2_17_pdst},
     {rob_uop_2_16_pdst},
     {rob_uop_2_15_pdst},
     {rob_uop_2_14_pdst},
     {rob_uop_2_13_pdst},
     {rob_uop_2_12_pdst},
     {rob_uop_2_11_pdst},
     {rob_uop_2_10_pdst},
     {rob_uop_2_9_pdst},
     {rob_uop_2_8_pdst},
     {rob_uop_2_7_pdst},
     {rob_uop_2_6_pdst},
     {rob_uop_2_5_pdst},
     {rob_uop_2_4_pdst},
     {rob_uop_2_3_pdst},
     {rob_uop_2_2_pdst},
     {rob_uop_2_1_pdst},
     {rob_uop_2_0_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0][6:0] _GEN_79 =
    {{rob_uop_2_31_stale_pdst},
     {rob_uop_2_30_stale_pdst},
     {rob_uop_2_29_stale_pdst},
     {rob_uop_2_28_stale_pdst},
     {rob_uop_2_27_stale_pdst},
     {rob_uop_2_26_stale_pdst},
     {rob_uop_2_25_stale_pdst},
     {rob_uop_2_24_stale_pdst},
     {rob_uop_2_23_stale_pdst},
     {rob_uop_2_22_stale_pdst},
     {rob_uop_2_21_stale_pdst},
     {rob_uop_2_20_stale_pdst},
     {rob_uop_2_19_stale_pdst},
     {rob_uop_2_18_stale_pdst},
     {rob_uop_2_17_stale_pdst},
     {rob_uop_2_16_stale_pdst},
     {rob_uop_2_15_stale_pdst},
     {rob_uop_2_14_stale_pdst},
     {rob_uop_2_13_stale_pdst},
     {rob_uop_2_12_stale_pdst},
     {rob_uop_2_11_stale_pdst},
     {rob_uop_2_10_stale_pdst},
     {rob_uop_2_9_stale_pdst},
     {rob_uop_2_8_stale_pdst},
     {rob_uop_2_7_stale_pdst},
     {rob_uop_2_6_stale_pdst},
     {rob_uop_2_5_stale_pdst},
     {rob_uop_2_4_stale_pdst},
     {rob_uop_2_3_stale_pdst},
     {rob_uop_2_2_stale_pdst},
     {rob_uop_2_1_stale_pdst},
     {rob_uop_2_0_stale_pdst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_80 =
    {{rob_uop_2_31_is_fencei},
     {rob_uop_2_30_is_fencei},
     {rob_uop_2_29_is_fencei},
     {rob_uop_2_28_is_fencei},
     {rob_uop_2_27_is_fencei},
     {rob_uop_2_26_is_fencei},
     {rob_uop_2_25_is_fencei},
     {rob_uop_2_24_is_fencei},
     {rob_uop_2_23_is_fencei},
     {rob_uop_2_22_is_fencei},
     {rob_uop_2_21_is_fencei},
     {rob_uop_2_20_is_fencei},
     {rob_uop_2_19_is_fencei},
     {rob_uop_2_18_is_fencei},
     {rob_uop_2_17_is_fencei},
     {rob_uop_2_16_is_fencei},
     {rob_uop_2_15_is_fencei},
     {rob_uop_2_14_is_fencei},
     {rob_uop_2_13_is_fencei},
     {rob_uop_2_12_is_fencei},
     {rob_uop_2_11_is_fencei},
     {rob_uop_2_10_is_fencei},
     {rob_uop_2_9_is_fencei},
     {rob_uop_2_8_is_fencei},
     {rob_uop_2_7_is_fencei},
     {rob_uop_2_6_is_fencei},
     {rob_uop_2_5_is_fencei},
     {rob_uop_2_4_is_fencei},
     {rob_uop_2_3_is_fencei},
     {rob_uop_2_2_is_fencei},
     {rob_uop_2_1_is_fencei},
     {rob_uop_2_0_is_fencei}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_81 =
    {{rob_uop_2_31_uses_ldq},
     {rob_uop_2_30_uses_ldq},
     {rob_uop_2_29_uses_ldq},
     {rob_uop_2_28_uses_ldq},
     {rob_uop_2_27_uses_ldq},
     {rob_uop_2_26_uses_ldq},
     {rob_uop_2_25_uses_ldq},
     {rob_uop_2_24_uses_ldq},
     {rob_uop_2_23_uses_ldq},
     {rob_uop_2_22_uses_ldq},
     {rob_uop_2_21_uses_ldq},
     {rob_uop_2_20_uses_ldq},
     {rob_uop_2_19_uses_ldq},
     {rob_uop_2_18_uses_ldq},
     {rob_uop_2_17_uses_ldq},
     {rob_uop_2_16_uses_ldq},
     {rob_uop_2_15_uses_ldq},
     {rob_uop_2_14_uses_ldq},
     {rob_uop_2_13_uses_ldq},
     {rob_uop_2_12_uses_ldq},
     {rob_uop_2_11_uses_ldq},
     {rob_uop_2_10_uses_ldq},
     {rob_uop_2_9_uses_ldq},
     {rob_uop_2_8_uses_ldq},
     {rob_uop_2_7_uses_ldq},
     {rob_uop_2_6_uses_ldq},
     {rob_uop_2_5_uses_ldq},
     {rob_uop_2_4_uses_ldq},
     {rob_uop_2_3_uses_ldq},
     {rob_uop_2_2_uses_ldq},
     {rob_uop_2_1_uses_ldq},
     {rob_uop_2_0_uses_ldq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_82 =
    {{rob_uop_2_31_uses_stq},
     {rob_uop_2_30_uses_stq},
     {rob_uop_2_29_uses_stq},
     {rob_uop_2_28_uses_stq},
     {rob_uop_2_27_uses_stq},
     {rob_uop_2_26_uses_stq},
     {rob_uop_2_25_uses_stq},
     {rob_uop_2_24_uses_stq},
     {rob_uop_2_23_uses_stq},
     {rob_uop_2_22_uses_stq},
     {rob_uop_2_21_uses_stq},
     {rob_uop_2_20_uses_stq},
     {rob_uop_2_19_uses_stq},
     {rob_uop_2_18_uses_stq},
     {rob_uop_2_17_uses_stq},
     {rob_uop_2_16_uses_stq},
     {rob_uop_2_15_uses_stq},
     {rob_uop_2_14_uses_stq},
     {rob_uop_2_13_uses_stq},
     {rob_uop_2_12_uses_stq},
     {rob_uop_2_11_uses_stq},
     {rob_uop_2_10_uses_stq},
     {rob_uop_2_9_uses_stq},
     {rob_uop_2_8_uses_stq},
     {rob_uop_2_7_uses_stq},
     {rob_uop_2_6_uses_stq},
     {rob_uop_2_5_uses_stq},
     {rob_uop_2_4_uses_stq},
     {rob_uop_2_3_uses_stq},
     {rob_uop_2_2_uses_stq},
     {rob_uop_2_1_uses_stq},
     {rob_uop_2_0_uses_stq}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_83 =
    {{rob_uop_2_31_is_sys_pc2epc},
     {rob_uop_2_30_is_sys_pc2epc},
     {rob_uop_2_29_is_sys_pc2epc},
     {rob_uop_2_28_is_sys_pc2epc},
     {rob_uop_2_27_is_sys_pc2epc},
     {rob_uop_2_26_is_sys_pc2epc},
     {rob_uop_2_25_is_sys_pc2epc},
     {rob_uop_2_24_is_sys_pc2epc},
     {rob_uop_2_23_is_sys_pc2epc},
     {rob_uop_2_22_is_sys_pc2epc},
     {rob_uop_2_21_is_sys_pc2epc},
     {rob_uop_2_20_is_sys_pc2epc},
     {rob_uop_2_19_is_sys_pc2epc},
     {rob_uop_2_18_is_sys_pc2epc},
     {rob_uop_2_17_is_sys_pc2epc},
     {rob_uop_2_16_is_sys_pc2epc},
     {rob_uop_2_15_is_sys_pc2epc},
     {rob_uop_2_14_is_sys_pc2epc},
     {rob_uop_2_13_is_sys_pc2epc},
     {rob_uop_2_12_is_sys_pc2epc},
     {rob_uop_2_11_is_sys_pc2epc},
     {rob_uop_2_10_is_sys_pc2epc},
     {rob_uop_2_9_is_sys_pc2epc},
     {rob_uop_2_8_is_sys_pc2epc},
     {rob_uop_2_7_is_sys_pc2epc},
     {rob_uop_2_6_is_sys_pc2epc},
     {rob_uop_2_5_is_sys_pc2epc},
     {rob_uop_2_4_is_sys_pc2epc},
     {rob_uop_2_3_is_sys_pc2epc},
     {rob_uop_2_2_is_sys_pc2epc},
     {rob_uop_2_1_is_sys_pc2epc},
     {rob_uop_2_0_is_sys_pc2epc}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_84 =
    {{rob_uop_2_31_flush_on_commit},
     {rob_uop_2_30_flush_on_commit},
     {rob_uop_2_29_flush_on_commit},
     {rob_uop_2_28_flush_on_commit},
     {rob_uop_2_27_flush_on_commit},
     {rob_uop_2_26_flush_on_commit},
     {rob_uop_2_25_flush_on_commit},
     {rob_uop_2_24_flush_on_commit},
     {rob_uop_2_23_flush_on_commit},
     {rob_uop_2_22_flush_on_commit},
     {rob_uop_2_21_flush_on_commit},
     {rob_uop_2_20_flush_on_commit},
     {rob_uop_2_19_flush_on_commit},
     {rob_uop_2_18_flush_on_commit},
     {rob_uop_2_17_flush_on_commit},
     {rob_uop_2_16_flush_on_commit},
     {rob_uop_2_15_flush_on_commit},
     {rob_uop_2_14_flush_on_commit},
     {rob_uop_2_13_flush_on_commit},
     {rob_uop_2_12_flush_on_commit},
     {rob_uop_2_11_flush_on_commit},
     {rob_uop_2_10_flush_on_commit},
     {rob_uop_2_9_flush_on_commit},
     {rob_uop_2_8_flush_on_commit},
     {rob_uop_2_7_flush_on_commit},
     {rob_uop_2_6_flush_on_commit},
     {rob_uop_2_5_flush_on_commit},
     {rob_uop_2_4_flush_on_commit},
     {rob_uop_2_3_flush_on_commit},
     {rob_uop_2_2_flush_on_commit},
     {rob_uop_2_1_flush_on_commit},
     {rob_uop_2_0_flush_on_commit}};	// rob.scala:310:28, :411:25
  wire [31:0][5:0] _GEN_85 =
    {{rob_uop_2_31_ldst},
     {rob_uop_2_30_ldst},
     {rob_uop_2_29_ldst},
     {rob_uop_2_28_ldst},
     {rob_uop_2_27_ldst},
     {rob_uop_2_26_ldst},
     {rob_uop_2_25_ldst},
     {rob_uop_2_24_ldst},
     {rob_uop_2_23_ldst},
     {rob_uop_2_22_ldst},
     {rob_uop_2_21_ldst},
     {rob_uop_2_20_ldst},
     {rob_uop_2_19_ldst},
     {rob_uop_2_18_ldst},
     {rob_uop_2_17_ldst},
     {rob_uop_2_16_ldst},
     {rob_uop_2_15_ldst},
     {rob_uop_2_14_ldst},
     {rob_uop_2_13_ldst},
     {rob_uop_2_12_ldst},
     {rob_uop_2_11_ldst},
     {rob_uop_2_10_ldst},
     {rob_uop_2_9_ldst},
     {rob_uop_2_8_ldst},
     {rob_uop_2_7_ldst},
     {rob_uop_2_6_ldst},
     {rob_uop_2_5_ldst},
     {rob_uop_2_4_ldst},
     {rob_uop_2_3_ldst},
     {rob_uop_2_2_ldst},
     {rob_uop_2_1_ldst},
     {rob_uop_2_0_ldst}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_86 =
    {{rob_uop_2_31_ldst_val},
     {rob_uop_2_30_ldst_val},
     {rob_uop_2_29_ldst_val},
     {rob_uop_2_28_ldst_val},
     {rob_uop_2_27_ldst_val},
     {rob_uop_2_26_ldst_val},
     {rob_uop_2_25_ldst_val},
     {rob_uop_2_24_ldst_val},
     {rob_uop_2_23_ldst_val},
     {rob_uop_2_22_ldst_val},
     {rob_uop_2_21_ldst_val},
     {rob_uop_2_20_ldst_val},
     {rob_uop_2_19_ldst_val},
     {rob_uop_2_18_ldst_val},
     {rob_uop_2_17_ldst_val},
     {rob_uop_2_16_ldst_val},
     {rob_uop_2_15_ldst_val},
     {rob_uop_2_14_ldst_val},
     {rob_uop_2_13_ldst_val},
     {rob_uop_2_12_ldst_val},
     {rob_uop_2_11_ldst_val},
     {rob_uop_2_10_ldst_val},
     {rob_uop_2_9_ldst_val},
     {rob_uop_2_8_ldst_val},
     {rob_uop_2_7_ldst_val},
     {rob_uop_2_6_ldst_val},
     {rob_uop_2_5_ldst_val},
     {rob_uop_2_4_ldst_val},
     {rob_uop_2_3_ldst_val},
     {rob_uop_2_2_ldst_val},
     {rob_uop_2_1_ldst_val},
     {rob_uop_2_0_ldst_val}};	// rob.scala:310:28, :411:25
  wire [31:0][1:0] _GEN_87 =
    {{rob_uop_2_31_dst_rtype},
     {rob_uop_2_30_dst_rtype},
     {rob_uop_2_29_dst_rtype},
     {rob_uop_2_28_dst_rtype},
     {rob_uop_2_27_dst_rtype},
     {rob_uop_2_26_dst_rtype},
     {rob_uop_2_25_dst_rtype},
     {rob_uop_2_24_dst_rtype},
     {rob_uop_2_23_dst_rtype},
     {rob_uop_2_22_dst_rtype},
     {rob_uop_2_21_dst_rtype},
     {rob_uop_2_20_dst_rtype},
     {rob_uop_2_19_dst_rtype},
     {rob_uop_2_18_dst_rtype},
     {rob_uop_2_17_dst_rtype},
     {rob_uop_2_16_dst_rtype},
     {rob_uop_2_15_dst_rtype},
     {rob_uop_2_14_dst_rtype},
     {rob_uop_2_13_dst_rtype},
     {rob_uop_2_12_dst_rtype},
     {rob_uop_2_11_dst_rtype},
     {rob_uop_2_10_dst_rtype},
     {rob_uop_2_9_dst_rtype},
     {rob_uop_2_8_dst_rtype},
     {rob_uop_2_7_dst_rtype},
     {rob_uop_2_6_dst_rtype},
     {rob_uop_2_5_dst_rtype},
     {rob_uop_2_4_dst_rtype},
     {rob_uop_2_3_dst_rtype},
     {rob_uop_2_2_dst_rtype},
     {rob_uop_2_1_dst_rtype},
     {rob_uop_2_0_dst_rtype}};	// rob.scala:310:28, :411:25
  wire [31:0]      _GEN_88 =
    {{rob_uop_2_31_fp_val},
     {rob_uop_2_30_fp_val},
     {rob_uop_2_29_fp_val},
     {rob_uop_2_28_fp_val},
     {rob_uop_2_27_fp_val},
     {rob_uop_2_26_fp_val},
     {rob_uop_2_25_fp_val},
     {rob_uop_2_24_fp_val},
     {rob_uop_2_23_fp_val},
     {rob_uop_2_22_fp_val},
     {rob_uop_2_21_fp_val},
     {rob_uop_2_20_fp_val},
     {rob_uop_2_19_fp_val},
     {rob_uop_2_18_fp_val},
     {rob_uop_2_17_fp_val},
     {rob_uop_2_16_fp_val},
     {rob_uop_2_15_fp_val},
     {rob_uop_2_14_fp_val},
     {rob_uop_2_13_fp_val},
     {rob_uop_2_12_fp_val},
     {rob_uop_2_11_fp_val},
     {rob_uop_2_10_fp_val},
     {rob_uop_2_9_fp_val},
     {rob_uop_2_8_fp_val},
     {rob_uop_2_7_fp_val},
     {rob_uop_2_6_fp_val},
     {rob_uop_2_5_fp_val},
     {rob_uop_2_4_fp_val},
     {rob_uop_2_3_fp_val},
     {rob_uop_2_2_fp_val},
     {rob_uop_2_1_fp_val},
     {rob_uop_2_0_fp_val}};	// rob.scala:310:28, :411:25
  wire             rbk_row_2 = _io_commit_rollback_T_2 & ~full;	// rob.scala:236:31, :425:{44,47}, :787:39
  wire             _io_commit_rbk_valids_2_output = rbk_row_2 & _GEN_59[com_idx];	// rob.scala:236:20, :324:31, :425:44, :427:40
  reg              block_commit_REG;	// rob.scala:540:94
  reg              block_commit_REG_1;	// rob.scala:540:131
  reg              block_commit_REG_2;	// rob.scala:540:123
  wire             block_commit =
    rob_state != 2'h1 & rob_state != 2'h3 | block_commit_REG | block_commit_REG_2;	// rob.scala:221:26, :419:36, :540:{33,47,61,94,113,123}
  assign will_commit_0 = can_commit_0 & ~can_throw_exception_0 & ~block_commit;	// rob.scala:398:49, :404:64, :540:113, :545:55, :547:{46,70}
  wire             _GEN_89 =
    rob_head_vals_0 & (~can_commit_0 | can_throw_exception_0) | block_commit;	// rob.scala:398:49, :404:64, :540:113, :548:46, :549:{29,44,72}
  assign will_commit_1 = can_commit_1 & ~can_throw_exception_1 & ~_GEN_89;	// rob.scala:398:49, :404:64, :545:55, :547:{46,70}, :549:72
  wire             _GEN_90 =
    rob_head_vals_1 & (~can_commit_1 | can_throw_exception_1) | _GEN_89;	// rob.scala:398:49, :404:64, :548:46, :549:{29,44,72}
  wire             exception_thrown =
    can_throw_exception_2 & ~_GEN_90 & ~will_commit_1 | can_throw_exception_1 & ~_GEN_89
    & ~will_commit_0 | can_throw_exception_0 & ~block_commit;	// rob.scala:398:49, :540:113, :545:{52,55,69,72,85}, :547:70, :549:72
  assign will_commit_2 =
    rob_head_vals_2 & ~_GEN_67[rob_head] & ~io_csr_stall & ~can_throw_exception_2
    & ~_GEN_90;	// rob.scala:224:29, :366:31, :398:49, :404:{43,67}, :545:55, :547:{46,70}, :549:72
  wire             _io_flush_bits_flush_typ_T = r_xcpt_uop_exc_cause != 64'h10;	// rob.scala:259:29, :556:50
  wire [4:0]       com_xcpt_uop_ftq_idx =
    rob_head_vals_0
      ? _GEN_15[com_idx]
      : rob_head_vals_1 ? _GEN_45[com_idx] : _GEN_75[com_idx];	// Mux.scala:47:69, rob.scala:236:20, :398:49, :411:25
  wire             com_xcpt_uop_edge_inst =
    rob_head_vals_0
      ? _GEN_16[com_idx]
      : rob_head_vals_1 ? _GEN_46[com_idx] : _GEN_76[com_idx];	// Mux.scala:47:69, rob.scala:236:20, :398:49, :411:25
  wire [5:0]       com_xcpt_uop_pc_lob =
    rob_head_vals_0
      ? _GEN_17[com_idx]
      : rob_head_vals_1 ? _GEN_47[com_idx] : _GEN_77[com_idx];	// Mux.scala:47:69, rob.scala:236:20, :398:49, :411:25
  wire             flush_commit_mask_0 = will_commit_0 & _GEN_24[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit_mask_1 = will_commit_1 & _GEN_54[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit_mask_2 = will_commit_2 & _GEN_84[com_idx];	// rob.scala:236:20, :411:25, :547:70, :571:75
  wire             flush_commit =
    flush_commit_mask_0 | flush_commit_mask_1 | flush_commit_mask_2;	// rob.scala:571:75, :572:48
  wire             _io_flush_valid_output = exception_thrown | flush_commit;	// rob.scala:545:85, :572:48, :573:36
  wire             _fflags_val_0_T = will_commit_0 & _GEN_28[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_0 = _fflags_val_0_T & ~_GEN_22[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  wire             _fflags_val_1_T = will_commit_1 & _GEN_58[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_1 = _fflags_val_1_T & ~_GEN_52[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  wire             _fflags_val_2_T = will_commit_2 & _GEN_88[com_idx];	// rob.scala:236:20, :411:25, :547:70, :601:27
  wire             fflags_val_2 = _fflags_val_2_T & ~_GEN_82[com_idx];	// rob.scala:236:20, :411:25, :601:27, :602:32, :603:7
  reg              r_partial_row;	// rob.scala:677:30
  wire             _empty_T = rob_head == rob_tail;	// rob.scala:224:29, :228:29, :686:33
  wire             finished_committing_row =
    (|{will_commit_2, will_commit_1, will_commit_0})
    & ({will_commit_2, will_commit_1, will_commit_0}
       ^ {rob_head_vals_2, rob_head_vals_1, rob_head_vals_0}) == 3'h0
    & ~(r_partial_row & _empty_T & ~maybe_full);	// rob.scala:239:29, :398:49, :547:70, :677:30, :684:{23,30}, :685:{19,26,42,50,59}, :686:{5,33,46,49}
  reg              pnr_maybe_at_tail;	// rob.scala:714:36
  wire             _io_ready_T = rob_state == 2'h1;	// rob.scala:221:26, :540:33, :716:33
  `ifndef SYNTHESIS	// rob.scala:333:14
    always @(posedge clock) begin	// rob.scala:333:14
      automatic logic [6:0] rob_pnr_idx;	// Cat.scala:30:58
      automatic logic       _GEN_91 = io_lxcpt_bits_cause != 5'h10;	// rob.scala:324:31, :392:33
      automatic logic       _GEN_92 =
        ~((will_commit_0 | will_commit_1 | will_commit_2)
          & (_io_commit_rbk_valids_0_output | _io_commit_rbk_valids_1_output
             | _io_commit_rbk_valids_2_output)) | reset;	// rob.scala:427:40, :430:{12,13,40,45,77}, :547:70
      automatic logic       _GEN_93;	// util.scala:363:52
      automatic logic [1:0] _GEN_94 =
        {1'h0, flush_commit_mask_0} + {1'h0, flush_commit_mask_1}
        + {1'h0, flush_commit_mask_2};	// Bitwise.scala:47:55, rob.scala:361:75, :370:59, :372:26, :571:75
      rob_pnr_idx = {rob_pnr, rob_pnr_lsb};	// Cat.scala:30:58, rob.scala:232:29, :233:29
      _GEN_93 = rob_pnr_idx < rob_head_idx;	// Cat.scala:30:58, util.scala:363:52
      if (io_enq_valids_0 & ~(~rob_tail_vals_0 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_0 & ~(io_enq_uops_0_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_6 & ~(_GEN[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_6 & ~(_GEN_7[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_8 & ~(_GEN[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_8 & ~(_GEN_7[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_9 & _GEN_91 & ~(_GEN_10[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_92) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_0 & ~_GEN[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_0 & ~_GEN_7[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_0 & _GEN_26[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_18[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_1 & ~_GEN[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_1 & ~_GEN_7[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_1 & _GEN_26[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_18[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_2 & ~_GEN[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_2 & ~_GEN_7[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_2 & _GEN_26[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_18[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_3 & ~_GEN[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_3 & ~_GEN_7[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_3 & _GEN_26[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_18[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_4 & ~_GEN[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_4 & ~_GEN_7[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_4 & _GEN_26[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_18[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_5 & ~_GEN[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_5 & ~_GEN_7[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_5 & _GEN_26[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_18[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (io_enq_valids_1 & ~(~rob_tail_vals_1 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_1 & ~(io_enq_uops_1_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_36 & ~(_GEN_29[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_36 & ~(_GEN_37[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_38 & ~(_GEN_29[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_38 & ~(_GEN_37[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_39 & _GEN_91 & ~(_GEN_40[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_92) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_30 & ~_GEN_29[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_30 & ~_GEN_37[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_30 & _GEN_56[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_48[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_31 & ~_GEN_29[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_31 & ~_GEN_37[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_31 & _GEN_56[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_48[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_32 & ~_GEN_29[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_32 & ~_GEN_37[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_32 & _GEN_56[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_48[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_33 & ~_GEN_29[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_33 & ~_GEN_37[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_33 & _GEN_56[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_48[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_34 & ~_GEN_29[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_34 & ~_GEN_37[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_34 & _GEN_56[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_48[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_35 & ~_GEN_29[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_35 & ~_GEN_37[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_35 & _GEN_56[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_48[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (io_enq_valids_2 & ~(~rob_tail_vals_2 | reset)) begin	// rob.scala:324:31, :333:{14,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:333:14
          $error("Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");	// rob.scala:333:14
        if (`STOP_COND_)	// rob.scala:333:14
          $fatal;	// rob.scala:333:14
      end
      if (io_enq_valids_2 & ~(io_enq_uops_2_rob_idx[6:2] == rob_tail | reset)) begin	// rob.scala:228:29, :334:{14,39,63}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:334:14
          $error("Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");	// rob.scala:334:14
        if (`STOP_COND_)	// rob.scala:334:14
          $fatal;	// rob.scala:334:14
      end
      if (_GEN_66 & ~(_GEN_59[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_66 & ~(_GEN_67[io_lsu_clr_bsy_0_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_68 & ~(_GEN_59[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :361:31, :365:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:365:16
          $error("Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");	// rob.scala:365:16
        if (`STOP_COND_)	// rob.scala:365:16
          $fatal;	// rob.scala:365:16
      end
      if (_GEN_68 & ~(_GEN_67[io_lsu_clr_bsy_1_bits[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :361:31, :366:{16,31}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:366:16
          $error("Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");	// rob.scala:366:16
        if (`STOP_COND_)	// rob.scala:366:16
          $fatal;	// rob.scala:366:16
      end
      if (_GEN_69 & _GEN_91 & ~(_GEN_70[io_lxcpt_bits_uop_rob_idx[6:2]] | reset)) begin	// rob.scala:236:31, :268:25, :390:26, :392:33, :394:15
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:394:15
          $error("Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");	// rob.scala:394:15
        if (`STOP_COND_)	// rob.scala:394:15
          $fatal;	// rob.scala:394:15
      end
      if (~_GEN_92) begin	// rob.scala:430:12
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:430:12
          $error("Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:430 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");	// rob.scala:430:12
        if (`STOP_COND_)	// rob.scala:430:12
          $fatal;	// rob.scala:430:12
      end
      if (~(~(_GEN_60 & ~_GEN_59[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_60 & ~_GEN_67[io_wb_resps_0_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_60 & _GEN_86[io_wb_resps_0_bits_uop_rob_idx[6:2]]
              & _GEN_78[io_wb_resps_0_bits_uop_rob_idx[6:2]] != io_wb_resps_0_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_61 & ~_GEN_59[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_61 & ~_GEN_67[io_wb_resps_1_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_61 & _GEN_86[io_wb_resps_1_bits_uop_rob_idx[6:2]]
              & _GEN_78[io_wb_resps_1_bits_uop_rob_idx[6:2]] != io_wb_resps_1_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_62 & ~_GEN_59[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_62 & ~_GEN_67[io_wb_resps_2_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_62 & _GEN_86[io_wb_resps_2_bits_uop_rob_idx[6:2]]
              & _GEN_78[io_wb_resps_2_bits_uop_rob_idx[6:2]] != io_wb_resps_2_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_63 & ~_GEN_59[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_63 & ~_GEN_67[io_wb_resps_3_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_63 & _GEN_86[io_wb_resps_3_bits_uop_rob_idx[6:2]]
              & _GEN_78[io_wb_resps_3_bits_uop_rob_idx[6:2]] != io_wb_resps_3_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_64 & ~_GEN_59[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_64 & ~_GEN_67[io_wb_resps_4_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_64 & _GEN_86[io_wb_resps_4_bits_uop_rob_idx[6:2]]
              & _GEN_78[io_wb_resps_4_bits_uop_rob_idx[6:2]] != io_wb_resps_4_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_65 & ~_GEN_59[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :324:31, :346:27, :514:{14,15,72}, :515:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:514:14
          $error("Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:514 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:514:14
        if (`STOP_COND_)	// rob.scala:514:14
          $fatal;	// rob.scala:514:14
      end
      if (~(~(_GEN_65 & ~_GEN_67[io_wb_resps_5_bits_uop_rob_idx[6:2]]) | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :366:31, :517:{14,15,72}, :518:16
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:517:14
          $error("Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:517 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:517:14
        if (`STOP_COND_)	// rob.scala:517:14
          $fatal;	// rob.scala:517:14
      end
      if (~(~(_GEN_65 & _GEN_86[io_wb_resps_5_bits_uop_rob_idx[6:2]]
              & _GEN_78[io_wb_resps_5_bits_uop_rob_idx[6:2]] != io_wb_resps_5_bits_uop_pdst)
            | reset)) begin	// rob.scala:236:31, :268:25, :346:27, :411:25, :520:{14,15,72}, :521:{34,51}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:520:14
          $error("Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:520 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");	// rob.scala:520:14
        if (`STOP_COND_)	// rob.scala:520:14
          $fatal;	// rob.scala:520:14
      end
      if (~(~(_GEN_94[1]) | reset)) begin	// Bitwise.scala:47:55, rob.scala:575:{9,10,40}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:575:9
          $error("Assertion failed: [rob] Can't commit multiple flush_on_commit instructions on one cycle\n    at rob.scala:575 assert(!(PopCount(flush_commit_mask) > 1.U),\n");	// rob.scala:575:9
        if (`STOP_COND_)	// rob.scala:575:9
          $fatal;	// rob.scala:575:9
      end
      if (~(~(will_commit_0 & ~_GEN_28[com_idx] & (|_rob_fflags_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_0_T & (_GEN_21[com_idx] | _GEN_22[com_idx])
              & (|_rob_fflags_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(will_commit_1 & ~_GEN_58[com_idx] & (|_rob_fflags_1_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_1_T & (_GEN_51[com_idx] | _GEN_52[com_idx])
              & (|_rob_fflags_1_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(will_commit_2 & ~_GEN_88[com_idx] & (|_rob_fflags_2_ext_R0_data))
            | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :547:70, :607:{12,13}, :608:{14,40}, :609:33
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:607:12
          $error("Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:607 assert (!(io.commit.valids(w) &&\n");	// rob.scala:607:12
        if (`STOP_COND_)	// rob.scala:607:12
          $fatal;	// rob.scala:607:12
      end
      if (~(~(_fflags_val_2_T & (_GEN_81[com_idx] | _GEN_82[com_idx])
              & (|_rob_fflags_2_ext_R0_data)) | reset)) begin	// rob.scala:236:20, :313:28, :411:25, :601:27, :609:33, :611:{12,13}, :613:{42,73}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:611:12
          $error("Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:611 assert (!(io.commit.valids(w) &&\n");	// rob.scala:611:12
        if (`STOP_COND_)	// rob.scala:611:12
          $fatal;	// rob.scala:611:12
      end
      if (~(~(exception_thrown & ~r_xcpt_val) | reset)) begin	// rob.scala:258:33, :545:85, :658:{10,11,30,33}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:658:10
          $error("Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:658 assert (!(exception_thrown && !r_xcpt_val),\n");	// rob.scala:658:10
        if (`STOP_COND_)	// rob.scala:658:10
          $fatal;	// rob.scala:658:10
      end
      if (~(~(empty & r_xcpt_val) | reset)) begin	// rob.scala:258:33, :661:{10,11,19}, :788:41
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:661:10
          $error("Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:661 assert (!(empty && r_xcpt_val),\n");	// rob.scala:661:10
        if (`STOP_COND_)	// rob.scala:661:10
          $fatal;	// rob.scala:661:10
      end
      if (~(~(exception_thrown & r_xcpt_uop_rob_idx[6:2] != rob_head) | reset)) begin	// rob.scala:224:29, :236:31, :259:29, :268:25, :545:85, :664:{10,11,34,68}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:664:10
          $error("Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:664 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n");	// rob.scala:664:10
        if (`STOP_COND_)	// rob.scala:664:10
          $fatal;	// rob.scala:664:10
      end
      if (~(_GEN_93 ^ rob_head_idx < rob_tail_idx ^ rob_pnr_idx >= rob_tail_idx
            | rob_pnr_idx == rob_tail_idx | reset)) begin	// Cat.scala:30:58, rob.scala:740:{9,10,75}, util.scala:363:{52,64,78}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:740:9
          $error("Assertion failed\n    at rob.scala:740 assert(!IsOlder(rob_pnr_idx, rob_head_idx, rob_tail_idx) || rob_pnr_idx === rob_tail_idx)\n");	// rob.scala:740:9
        if (`STOP_COND_)	// rob.scala:740:9
          $fatal;	// rob.scala:740:9
      end
      if (~(rob_tail_idx < rob_head_idx ^ _GEN_93 ^ rob_tail_idx >= rob_pnr_idx | full
            | reset)) begin	// Cat.scala:30:58, rob.scala:743:{9,10}, :787:39, util.scala:363:{52,64}
        if (`ASSERT_VERBOSE_COND_)	// rob.scala:743:9
          $error("Assertion failed\n    at rob.scala:743 assert(!IsOlder(rob_tail_idx, rob_pnr_idx, rob_head_idx) || full)\n");	// rob.scala:743:9
        if (`STOP_COND_)	// rob.scala:743:9
          $fatal;	// rob.scala:743:9
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire             _GEN_95 =
    _io_commit_rollback_T_2 & (rob_tail != rob_head | maybe_full);	// rob.scala:224:29, :228:29, :236:31, :239:29, :750:{34,47,60}
  wire             rob_deq = _GEN_95 | finished_committing_row;	// rob.scala:685:59, :688:34, :750:{34,76}, :754:13
  assign full = rob_tail == rob_head & maybe_full;	// rob.scala:224:29, :228:29, :239:29, :787:{26,39}
  assign empty = _empty_T & {rob_head_vals_2, rob_head_vals_1, rob_head_vals_0} == 3'h0;	// rob.scala:398:49, :686:33, :788:{41,59,66}
  reg              REG;	// rob.scala:808:30
  reg              REG_1;	// rob.scala:808:22
  reg              REG_2;	// rob.scala:824:22
  reg              io_com_load_is_at_rob_head_REG;	// rob.scala:865:40
  always @(posedge clock) begin
    automatic logic             _GEN_96;	// rob.scala:324:31
    automatic logic             _GEN_97;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_98;	// rob.scala:324:31
    automatic logic             _GEN_99;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_100;	// rob.scala:324:31
    automatic logic             _GEN_101;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_102;	// rob.scala:324:31
    automatic logic             _GEN_103;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_104;	// rob.scala:324:31
    automatic logic             _GEN_105;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_106;	// rob.scala:324:31
    automatic logic             _GEN_107;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_108;	// rob.scala:324:31
    automatic logic             _GEN_109;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_110;	// rob.scala:324:31
    automatic logic             _GEN_111;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_112;	// rob.scala:324:31
    automatic logic             _GEN_113;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_114;	// rob.scala:324:31
    automatic logic             _GEN_115;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_116;	// rob.scala:324:31
    automatic logic             _GEN_117;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_118;	// rob.scala:324:31
    automatic logic             _GEN_119;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_120;	// rob.scala:324:31
    automatic logic             _GEN_121;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_122;	// rob.scala:324:31
    automatic logic             _GEN_123;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_124;	// rob.scala:324:31
    automatic logic             _GEN_125;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_126;	// rob.scala:324:31
    automatic logic             _GEN_127;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_128;	// rob.scala:324:31
    automatic logic             _GEN_129;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_130;	// rob.scala:324:31
    automatic logic             _GEN_131;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_132;	// rob.scala:324:31
    automatic logic             _GEN_133;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_134;	// rob.scala:324:31
    automatic logic             _GEN_135;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_136;	// rob.scala:324:31
    automatic logic             _GEN_137;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_138;	// rob.scala:324:31
    automatic logic             _GEN_139;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_140;	// rob.scala:324:31
    automatic logic             _GEN_141;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_142;	// rob.scala:324:31
    automatic logic             _GEN_143;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_144;	// rob.scala:324:31
    automatic logic             _GEN_145;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_146;	// rob.scala:324:31
    automatic logic             _GEN_147;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_148;	// rob.scala:324:31
    automatic logic             _GEN_149;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_150;	// rob.scala:324:31
    automatic logic             _GEN_151;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_152;	// rob.scala:324:31
    automatic logic             _GEN_153;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_154;	// rob.scala:324:31
    automatic logic             _GEN_155;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_156;	// rob.scala:324:31
    automatic logic             _GEN_157;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_158;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T =
      io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_159;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_160;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_161;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_162;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_163;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_164;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_165;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_166;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_167;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_168;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_169;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_170;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_171;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_172;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_173;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_174;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_175;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_176;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_177;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_178;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_179;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_180;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_181;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_182;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_183;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_184;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_185;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_186;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_187;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_188;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_189;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_190;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_4 =
      io_enq_uops_0_uses_ldq | io_enq_uops_0_uses_stq & ~io_enq_uops_0_is_fence
      | io_enq_uops_0_is_br | io_enq_uops_0_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_191;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_192;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_193;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_194;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_195;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_196;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_197;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_198;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_199;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_200;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_201;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_202;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_203;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_204;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_205;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_206;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_207;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_208;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_209;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_210;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_211;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_212;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_213;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_214;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_215;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_216;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_217;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_218;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_219;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_220;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_221;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_222;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_223 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :347:31
    automatic logic             _GEN_224 = _GEN_0 & _GEN_223;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_225 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_226 = _GEN_0 & _GEN_225;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_227 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_228 = _GEN_0 & _GEN_227;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_229 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_230 = _GEN_0 & _GEN_229;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_231 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_232 = _GEN_0 & _GEN_231;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_233 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_234 = _GEN_0 & _GEN_233;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_235 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_236 = _GEN_0 & _GEN_235;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_237 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_238 = _GEN_0 & _GEN_237;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_239 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_240 = _GEN_0 & _GEN_239;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_241 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_242 = _GEN_0 & _GEN_241;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_243 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_244 = _GEN_0 & _GEN_243;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_245 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_246 = _GEN_0 & _GEN_245;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_247 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_248 = _GEN_0 & _GEN_247;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_249 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_250 = _GEN_0 & _GEN_249;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_251 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_252 = _GEN_0 & _GEN_251;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_253 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_254 = _GEN_0 & _GEN_253;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_255 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_256 = _GEN_0 & _GEN_255;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_257 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_258 = _GEN_0 & _GEN_257;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_259 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_260 = _GEN_0 & _GEN_259;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_261 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_262 = _GEN_0 & _GEN_261;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_263 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_264 = _GEN_0 & _GEN_263;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_265 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_266 = _GEN_0 & _GEN_265;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_267 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_268 = _GEN_0 & _GEN_267;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_269 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_270 = _GEN_0 & _GEN_269;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_271 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_272 = _GEN_0 & _GEN_271;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_273 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_274 = _GEN_0 & _GEN_273;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_275 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_276 = _GEN_0 & _GEN_275;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_277 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_278 = _GEN_0 & _GEN_277;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_279 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_280 = _GEN_0 & _GEN_279;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_281 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_282 = _GEN_0 & _GEN_281;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_283 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_284 = _GEN_0 & _GEN_283;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_285 =
      _GEN_0 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_286 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :347:31
    automatic logic             _GEN_287 = _GEN_286 | _GEN_224;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_288;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_289 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_290 = _GEN_289 | _GEN_226;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_291;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_292 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_293 = _GEN_292 | _GEN_228;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_294;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_295 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_296 = _GEN_295 | _GEN_230;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_297;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_298 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_299 = _GEN_298 | _GEN_232;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_300;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_301 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_302 = _GEN_301 | _GEN_234;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_303;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_304 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_305 = _GEN_304 | _GEN_236;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_306;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_307 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_308 = _GEN_307 | _GEN_238;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_309;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_310 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_311 = _GEN_310 | _GEN_240;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_312;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_313 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_314 = _GEN_313 | _GEN_242;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_315;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_316 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_317 = _GEN_316 | _GEN_244;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_318;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_319 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_320 = _GEN_319 | _GEN_246;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_321;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_322 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_323 = _GEN_322 | _GEN_248;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_324;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_325 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_326 = _GEN_325 | _GEN_250;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_327;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_328 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_329 = _GEN_328 | _GEN_252;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_330;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_331 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_332 = _GEN_331 | _GEN_254;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_333;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_334 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_335 = _GEN_334 | _GEN_256;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_336;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_337 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_338 = _GEN_337 | _GEN_258;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_339;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_340 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_341 = _GEN_340 | _GEN_260;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_342;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_343 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_344 = _GEN_343 | _GEN_262;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_345;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_346 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_347 = _GEN_346 | _GEN_264;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_348;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_349 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_350 = _GEN_349 | _GEN_266;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_351;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_352 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_353 = _GEN_352 | _GEN_268;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_354;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_355 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_356 = _GEN_355 | _GEN_270;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_357;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_358 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_359 = _GEN_358 | _GEN_272;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_360;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_361 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_362 = _GEN_361 | _GEN_274;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_363;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_364 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_365 = _GEN_364 | _GEN_276;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_366;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_367 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_368 = _GEN_367 | _GEN_278;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_369;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_370 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_371 = _GEN_370 | _GEN_280;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_372;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_373 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_374 = _GEN_373 | _GEN_282;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_375;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_376 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_377 = _GEN_376 | _GEN_284;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_378;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_379 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_285;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_380;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_381;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_382;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_383;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_384;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_385;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_386;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_387;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_388;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_389;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_390;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_391;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_392;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_393;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_394;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_395;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_396;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_397;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_398;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_399;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_400;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_401;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_402;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_403;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_404;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_405;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_406;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_407;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_408;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_409;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_410;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_411;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_412;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_413 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :347:31
    automatic logic             _GEN_414 = _GEN_2 & _GEN_413;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_415 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_416 = _GEN_2 & _GEN_415;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_417 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_418 = _GEN_2 & _GEN_417;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_419 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_420 = _GEN_2 & _GEN_419;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_421 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_422 = _GEN_2 & _GEN_421;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_423 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_424 = _GEN_2 & _GEN_423;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_425 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_426 = _GEN_2 & _GEN_425;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_427 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_428 = _GEN_2 & _GEN_427;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_429 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_430 = _GEN_2 & _GEN_429;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_431 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_432 = _GEN_2 & _GEN_431;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_433 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_434 = _GEN_2 & _GEN_433;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_435 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_436 = _GEN_2 & _GEN_435;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_437 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_438 = _GEN_2 & _GEN_437;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_439 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_440 = _GEN_2 & _GEN_439;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_441 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_442 = _GEN_2 & _GEN_441;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_443 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_444 = _GEN_2 & _GEN_443;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_445 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_446 = _GEN_2 & _GEN_445;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_447 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_448 = _GEN_2 & _GEN_447;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_449 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_450 = _GEN_2 & _GEN_449;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_451 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_452 = _GEN_2 & _GEN_451;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_453 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_454 = _GEN_2 & _GEN_453;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_455 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_456 = _GEN_2 & _GEN_455;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_457 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_458 = _GEN_2 & _GEN_457;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_459 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_460 = _GEN_2 & _GEN_459;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_461 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_462 = _GEN_2 & _GEN_461;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_463 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_464 = _GEN_2 & _GEN_463;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_465 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_466 = _GEN_2 & _GEN_465;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_467 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_468 = _GEN_2 & _GEN_467;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_469 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_470 = _GEN_2 & _GEN_469;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_471 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_472 = _GEN_2 & _GEN_471;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_473 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_474 = _GEN_2 & _GEN_473;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_475 =
      _GEN_2 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_476 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :347:31
    automatic logic             _GEN_477 = _GEN_476 | _GEN_414;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_478;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_479 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_480 = _GEN_479 | _GEN_416;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_481;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_482 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_483 = _GEN_482 | _GEN_418;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_484;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_485 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_486 = _GEN_485 | _GEN_420;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_487;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_488 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_489 = _GEN_488 | _GEN_422;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_490;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_491 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_492 = _GEN_491 | _GEN_424;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_493;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_494 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_495 = _GEN_494 | _GEN_426;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_496;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_497 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_498 = _GEN_497 | _GEN_428;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_499;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_500 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_501 = _GEN_500 | _GEN_430;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_502;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_503 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_504 = _GEN_503 | _GEN_432;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_505;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_506 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_507 = _GEN_506 | _GEN_434;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_508;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_509 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_510 = _GEN_509 | _GEN_436;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_511;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_512 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_513 = _GEN_512 | _GEN_438;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_514;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_515 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_516 = _GEN_515 | _GEN_440;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_517;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_518 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_519 = _GEN_518 | _GEN_442;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_520;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_521 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_522 = _GEN_521 | _GEN_444;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_523;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_524 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_525 = _GEN_524 | _GEN_446;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_526;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_527 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_528 = _GEN_527 | _GEN_448;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_529;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_530 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_531 = _GEN_530 | _GEN_450;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_532;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_533 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_534 = _GEN_533 | _GEN_452;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_535;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_536 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_537 = _GEN_536 | _GEN_454;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_538;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_539 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_540 = _GEN_539 | _GEN_456;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_541;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_542 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_543 = _GEN_542 | _GEN_458;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_544;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_545 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_546 = _GEN_545 | _GEN_460;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_547;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_548 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_549 = _GEN_548 | _GEN_462;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_550;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_551 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_552 = _GEN_551 | _GEN_464;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_553;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_554 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_555 = _GEN_554 | _GEN_466;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_556;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_557 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_558 = _GEN_557 | _GEN_468;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_559;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_560 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_561 = _GEN_560 | _GEN_470;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_562;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_563 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_564 = _GEN_563 | _GEN_472;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_565;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_566 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_567 = _GEN_566 | _GEN_474;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_568;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_569 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_475;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_570;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_571;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_572;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_573;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_574;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_575;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_576;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_577;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_578;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_579;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_580;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_581;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_582;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_583;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_584;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_585;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_586;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_587;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_588;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_589;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_590;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_591;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_592;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_593;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_594;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_595;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_596;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_597;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_598;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_599;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_600;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_601;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_602;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_603 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :347:31
    automatic logic             _GEN_604 = _GEN_4 & _GEN_603;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_605 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_606 = _GEN_4 & _GEN_605;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_607 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_608 = _GEN_4 & _GEN_607;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_609 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_610 = _GEN_4 & _GEN_609;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_611 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_612 = _GEN_4 & _GEN_611;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_613 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_614 = _GEN_4 & _GEN_613;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_615 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_616 = _GEN_4 & _GEN_615;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_617 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_618 = _GEN_4 & _GEN_617;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_619 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_620 = _GEN_4 & _GEN_619;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_621 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_622 = _GEN_4 & _GEN_621;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_623 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_624 = _GEN_4 & _GEN_623;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_625 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_626 = _GEN_4 & _GEN_625;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_627 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_628 = _GEN_4 & _GEN_627;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_629 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_630 = _GEN_4 & _GEN_629;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_631 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_632 = _GEN_4 & _GEN_631;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_633 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_634 = _GEN_4 & _GEN_633;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_635 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_636 = _GEN_4 & _GEN_635;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_637 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_638 = _GEN_4 & _GEN_637;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_639 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_640 = _GEN_4 & _GEN_639;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_641 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_642 = _GEN_4 & _GEN_641;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_643 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_644 = _GEN_4 & _GEN_643;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_645 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_646 = _GEN_4 & _GEN_645;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_647 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_648 = _GEN_4 & _GEN_647;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_649 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_650 = _GEN_4 & _GEN_649;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_651 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_652 = _GEN_4 & _GEN_651;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_653 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_654 = _GEN_4 & _GEN_653;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_655 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_656 = _GEN_4 & _GEN_655;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_657 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_658 = _GEN_4 & _GEN_657;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_659 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_660 = _GEN_4 & _GEN_659;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_661 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_662 = _GEN_4 & _GEN_661;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_663 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_664 = _GEN_4 & _GEN_663;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_665 =
      _GEN_4 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_666 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :347:31
    automatic logic             _GEN_667 = _GEN_666 | _GEN_604;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_668;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_669 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_670 = _GEN_669 | _GEN_606;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_671;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_672 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_673 = _GEN_672 | _GEN_608;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_674;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_675 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_676 = _GEN_675 | _GEN_610;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_677;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_678 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_679 = _GEN_678 | _GEN_612;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_680;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_681 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_682 = _GEN_681 | _GEN_614;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_683;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_684 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_685 = _GEN_684 | _GEN_616;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_686;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_687 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_688 = _GEN_687 | _GEN_618;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_689;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_690 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_691 = _GEN_690 | _GEN_620;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_692;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_693 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_694 = _GEN_693 | _GEN_622;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_695;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_696 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_697 = _GEN_696 | _GEN_624;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_698;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_699 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_700 = _GEN_699 | _GEN_626;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_701;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_702 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_703 = _GEN_702 | _GEN_628;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_704;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_705 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_706 = _GEN_705 | _GEN_630;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_707;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_708 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_709 = _GEN_708 | _GEN_632;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_710;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_711 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_712 = _GEN_711 | _GEN_634;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_713;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_714 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_715 = _GEN_714 | _GEN_636;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_716;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_717 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_718 = _GEN_717 | _GEN_638;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_719;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_720 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_721 = _GEN_720 | _GEN_640;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_722;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_723 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_724 = _GEN_723 | _GEN_642;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_725;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_726 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_727 = _GEN_726 | _GEN_644;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_728;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_729 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_730 = _GEN_729 | _GEN_646;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_731;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_732 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_733 = _GEN_732 | _GEN_648;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_734;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_735 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_736 = _GEN_735 | _GEN_650;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_737;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_738 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_739 = _GEN_738 | _GEN_652;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_740;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_741 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_742 = _GEN_741 | _GEN_654;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_743;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_744 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_745 = _GEN_744 | _GEN_656;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_746;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_747 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_748 = _GEN_747 | _GEN_658;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_749;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_750 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_751 = _GEN_750 | _GEN_660;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_752;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_753 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_754 = _GEN_753 | _GEN_662;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_755;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_756 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :347:31
    automatic logic             _GEN_757 = _GEN_756 | _GEN_664;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_758;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_759 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_665;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_760;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_761;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_762;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_763;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_764;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_765;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_766;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_767;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_768;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_769;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_770;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_771;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_772;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_773;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_774;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_775;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_776;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_777;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_778;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_779;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_780;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_781;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_782;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_783;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_784;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_785;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_786;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_787;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_788;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_789;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_790;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_791;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_792;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_793 = io_lsu_clr_bsy_0_bits[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :363:26
    automatic logic             _GEN_794;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_795 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_796;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_797 = io_lsu_clr_bsy_0_bits[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_798;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_799 = io_lsu_clr_bsy_0_bits[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_800;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_801 = io_lsu_clr_bsy_0_bits[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_802;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_803 = io_lsu_clr_bsy_0_bits[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_804;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_805 = io_lsu_clr_bsy_0_bits[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_806;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_807 = io_lsu_clr_bsy_0_bits[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_808;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_809 = io_lsu_clr_bsy_0_bits[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_810;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_811 = io_lsu_clr_bsy_0_bits[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_812;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_813 = io_lsu_clr_bsy_0_bits[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_814;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_815 = io_lsu_clr_bsy_0_bits[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_816;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_817 = io_lsu_clr_bsy_0_bits[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_818;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_819 = io_lsu_clr_bsy_0_bits[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_820;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_821 = io_lsu_clr_bsy_0_bits[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_822;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_823 = io_lsu_clr_bsy_0_bits[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_824;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_825 = io_lsu_clr_bsy_0_bits[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_826;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_827 = io_lsu_clr_bsy_0_bits[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_828;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_829 = io_lsu_clr_bsy_0_bits[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_830;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_831 = io_lsu_clr_bsy_0_bits[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_832;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_833 = io_lsu_clr_bsy_0_bits[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_834;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_835 = io_lsu_clr_bsy_0_bits[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_836;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_837 = io_lsu_clr_bsy_0_bits[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_838;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_839 = io_lsu_clr_bsy_0_bits[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_840;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_841 = io_lsu_clr_bsy_0_bits[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_842;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_843 = io_lsu_clr_bsy_0_bits[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_844;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_845 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_846;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_847 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_848;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_849 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_850;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_851 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_852;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_853 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :363:26
    automatic logic             _GEN_854;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_855;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_856;	// rob.scala:363:26
    automatic logic             _GEN_857;	// rob.scala:363:26
    automatic logic             _GEN_858;	// rob.scala:363:26
    automatic logic             _GEN_859;	// rob.scala:363:26
    automatic logic             _GEN_860;	// rob.scala:363:26
    automatic logic             _GEN_861;	// rob.scala:363:26
    automatic logic             _GEN_862;	// rob.scala:363:26
    automatic logic             _GEN_863;	// rob.scala:363:26
    automatic logic             _GEN_864;	// rob.scala:363:26
    automatic logic             _GEN_865;	// rob.scala:363:26
    automatic logic             _GEN_866;	// rob.scala:363:26
    automatic logic             _GEN_867;	// rob.scala:363:26
    automatic logic             _GEN_868;	// rob.scala:363:26
    automatic logic             _GEN_869;	// rob.scala:363:26
    automatic logic             _GEN_870;	// rob.scala:363:26
    automatic logic             _GEN_871;	// rob.scala:363:26
    automatic logic             _GEN_872;	// rob.scala:363:26
    automatic logic             _GEN_873;	// rob.scala:363:26
    automatic logic             _GEN_874;	// rob.scala:363:26
    automatic logic             _GEN_875;	// rob.scala:363:26
    automatic logic             _GEN_876;	// rob.scala:363:26
    automatic logic             _GEN_877;	// rob.scala:363:26
    automatic logic             _GEN_878;	// rob.scala:363:26
    automatic logic             _GEN_879;	// rob.scala:363:26
    automatic logic             _GEN_880;	// rob.scala:363:26
    automatic logic             _GEN_881;	// rob.scala:363:26
    automatic logic             _GEN_882;	// rob.scala:363:26
    automatic logic             _GEN_883;	// rob.scala:363:26
    automatic logic             _GEN_884;	// rob.scala:363:26
    automatic logic             _GEN_885;	// rob.scala:363:26
    automatic logic             _GEN_886;	// rob.scala:363:26
    automatic logic             _GEN_887 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :391:59
    automatic logic             _GEN_888 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_889 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_890 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_891 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_892 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_893 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_894 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_895 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_896 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_897 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_898 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_899 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_900 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_901 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_902 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_903 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_904 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_905 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_906 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_907 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_908 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_909 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_910 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_911 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_912 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_913 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_914 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_915 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_916 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_917 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :391:59
    automatic logic             _GEN_918 = com_idx == 5'h0;	// rob.scala:224:29, :236:20, :434:30
    automatic logic             _GEN_919;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_920 = com_idx == 5'h1;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_921;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_922 = com_idx == 5'h2;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_923;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_924 = com_idx == 5'h3;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_925;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_926 = com_idx == 5'h4;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_927;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_928 = com_idx == 5'h5;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_929;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_930 = com_idx == 5'h6;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_931;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_932 = com_idx == 5'h7;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_933;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_934 = com_idx == 5'h8;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_935;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_936 = com_idx == 5'h9;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_937;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_938 = com_idx == 5'hA;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_939;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_940 = com_idx == 5'hB;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_941;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_942 = com_idx == 5'hC;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_943;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_944 = com_idx == 5'hD;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_945;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_946 = com_idx == 5'hE;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_947;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_948 = com_idx == 5'hF;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_949;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_950 = com_idx == 5'h10;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_951;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_952 = com_idx == 5'h11;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_953;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_954 = com_idx == 5'h12;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_955;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_956 = com_idx == 5'h13;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_957;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_958 = com_idx == 5'h14;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_959;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_960 = com_idx == 5'h15;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_961;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_962 = com_idx == 5'h16;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_963;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_964 = com_idx == 5'h17;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_965;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_966 = com_idx == 5'h18;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_967;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_968 = com_idx == 5'h19;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_969;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_970 = com_idx == 5'h1A;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_971;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_972 = com_idx == 5'h1B;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_973;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_974 = com_idx == 5'h1C;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_975;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_976 = com_idx == 5'h1D;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_977;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_978 = com_idx == 5'h1E;	// rob.scala:236:20, :324:31, :434:30
    automatic logic             _GEN_979;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_980;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [15:0]      _GEN_981;	// util.scala:118:51
    automatic logic [15:0]      _GEN_982;	// util.scala:118:51
    automatic logic [15:0]      _GEN_983;	// util.scala:118:51
    automatic logic [15:0]      _GEN_984;	// util.scala:118:51
    automatic logic [15:0]      _GEN_985;	// util.scala:118:51
    automatic logic [15:0]      _GEN_986;	// util.scala:118:51
    automatic logic [15:0]      _GEN_987;	// util.scala:118:51
    automatic logic [15:0]      _GEN_988;	// util.scala:118:51
    automatic logic [15:0]      _GEN_989;	// util.scala:118:51
    automatic logic [15:0]      _GEN_990;	// util.scala:118:51
    automatic logic [15:0]      _GEN_991;	// util.scala:118:51
    automatic logic [15:0]      _GEN_992;	// util.scala:118:51
    automatic logic [15:0]      _GEN_993;	// util.scala:118:51
    automatic logic [15:0]      _GEN_994;	// util.scala:118:51
    automatic logic [15:0]      _GEN_995;	// util.scala:118:51
    automatic logic [15:0]      _GEN_996;	// util.scala:118:51
    automatic logic [15:0]      _GEN_997;	// util.scala:118:51
    automatic logic [15:0]      _GEN_998;	// util.scala:118:51
    automatic logic [15:0]      _GEN_999;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1000;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1001;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1002;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1003;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1004;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1005;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1006;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1007;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1008;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1009;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1010;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1011;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1012;	// util.scala:118:51
    automatic logic             rob_head_uses_ldq_0;	// rob.scala:484:26
    automatic logic             _GEN_1013;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1014;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1015;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1016;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1017;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1018;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1019;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1020;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1021;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1022;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1023;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1024;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1025;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1026;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1027;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1028;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1029;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1030;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1031;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1032;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1033;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1034;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1035;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1036;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1037;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1038;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1039;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1040;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1041;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1042;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1043;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1044;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T_2 =
      io_enq_uops_1_is_fence | io_enq_uops_1_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_1045;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1046;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1047;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1048;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1049;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1050;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1051;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1052;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1053;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1054;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1055;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1056;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1057;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1058;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1059;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1060;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1061;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1062;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1063;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1064;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1065;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1066;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1067;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1068;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1069;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1070;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1071;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1072;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1073;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1074;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1075;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1076;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_9 =
      io_enq_uops_1_uses_ldq | io_enq_uops_1_uses_stq & ~io_enq_uops_1_is_fence
      | io_enq_uops_1_is_br | io_enq_uops_1_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_1077;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1078;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1079;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1080;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1081;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1082;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1083;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1084;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1085;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1086;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1087;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1088;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1089;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1090;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1091;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1092;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1093;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1094;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1095;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1096;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1097;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1098;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1099;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1100;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1101;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1102;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1103;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1104;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1105;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1106;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1107;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1108;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1109 = _GEN_30 & _GEN_223;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1110 = _GEN_30 & _GEN_225;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1111 = _GEN_30 & _GEN_227;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1112 = _GEN_30 & _GEN_229;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1113 = _GEN_30 & _GEN_231;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1114 = _GEN_30 & _GEN_233;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1115 = _GEN_30 & _GEN_235;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1116 = _GEN_30 & _GEN_237;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1117 = _GEN_30 & _GEN_239;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1118 = _GEN_30 & _GEN_241;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1119 = _GEN_30 & _GEN_243;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1120 = _GEN_30 & _GEN_245;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1121 = _GEN_30 & _GEN_247;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1122 = _GEN_30 & _GEN_249;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1123 = _GEN_30 & _GEN_251;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1124 = _GEN_30 & _GEN_253;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1125 = _GEN_30 & _GEN_255;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1126 = _GEN_30 & _GEN_257;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1127 = _GEN_30 & _GEN_259;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1128 = _GEN_30 & _GEN_261;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1129 = _GEN_30 & _GEN_263;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1130 = _GEN_30 & _GEN_265;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1131 = _GEN_30 & _GEN_267;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1132 = _GEN_30 & _GEN_269;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1133 = _GEN_30 & _GEN_271;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1134 = _GEN_30 & _GEN_273;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1135 = _GEN_30 & _GEN_275;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1136 = _GEN_30 & _GEN_277;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1137 = _GEN_30 & _GEN_279;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1138 = _GEN_30 & _GEN_281;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1139 = _GEN_30 & _GEN_283;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1140 =
      _GEN_30 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1141 = _GEN_286 | _GEN_1109;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1142;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1143 = _GEN_289 | _GEN_1110;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1144;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1145 = _GEN_292 | _GEN_1111;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1146;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1147 = _GEN_295 | _GEN_1112;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1148;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1149 = _GEN_298 | _GEN_1113;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1150;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1151 = _GEN_301 | _GEN_1114;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1152;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1153 = _GEN_304 | _GEN_1115;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1154;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1155 = _GEN_307 | _GEN_1116;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1156;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1157 = _GEN_310 | _GEN_1117;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1158;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1159 = _GEN_313 | _GEN_1118;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1160;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1161 = _GEN_316 | _GEN_1119;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1162;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1163 = _GEN_319 | _GEN_1120;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1164;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1165 = _GEN_322 | _GEN_1121;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1166;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1167 = _GEN_325 | _GEN_1122;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1168;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1169 = _GEN_328 | _GEN_1123;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1170;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1171 = _GEN_331 | _GEN_1124;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1172;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1173 = _GEN_334 | _GEN_1125;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1174;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1175 = _GEN_337 | _GEN_1126;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1176;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1177 = _GEN_340 | _GEN_1127;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1178;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1179 = _GEN_343 | _GEN_1128;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1180;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1181 = _GEN_346 | _GEN_1129;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1182;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1183 = _GEN_349 | _GEN_1130;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1184;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1185 = _GEN_352 | _GEN_1131;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1186;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1187 = _GEN_355 | _GEN_1132;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1188;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1189 = _GEN_358 | _GEN_1133;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1190;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1191 = _GEN_361 | _GEN_1134;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1192;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1193 = _GEN_364 | _GEN_1135;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1194;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1195 = _GEN_367 | _GEN_1136;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1196;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1197 = _GEN_370 | _GEN_1137;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1198;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1199 = _GEN_373 | _GEN_1138;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1200;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1201 = _GEN_376 | _GEN_1139;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1202;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1203 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_1140;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_1204;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1205;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1206;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1207;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1208;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1209;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1210;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1211;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1212;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1213;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1214;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1215;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1216;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1217;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1218;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1219;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1220;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1221;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1222;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1223;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1224;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1225;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1226;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1227;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1228;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1229;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1230;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1231;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1232;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1233;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1234;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1235;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1236;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1237 = _GEN_32 & _GEN_413;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1238 = _GEN_32 & _GEN_415;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1239 = _GEN_32 & _GEN_417;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1240 = _GEN_32 & _GEN_419;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1241 = _GEN_32 & _GEN_421;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1242 = _GEN_32 & _GEN_423;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1243 = _GEN_32 & _GEN_425;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1244 = _GEN_32 & _GEN_427;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1245 = _GEN_32 & _GEN_429;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1246 = _GEN_32 & _GEN_431;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1247 = _GEN_32 & _GEN_433;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1248 = _GEN_32 & _GEN_435;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1249 = _GEN_32 & _GEN_437;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1250 = _GEN_32 & _GEN_439;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1251 = _GEN_32 & _GEN_441;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1252 = _GEN_32 & _GEN_443;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1253 = _GEN_32 & _GEN_445;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1254 = _GEN_32 & _GEN_447;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1255 = _GEN_32 & _GEN_449;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1256 = _GEN_32 & _GEN_451;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1257 = _GEN_32 & _GEN_453;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1258 = _GEN_32 & _GEN_455;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1259 = _GEN_32 & _GEN_457;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1260 = _GEN_32 & _GEN_459;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1261 = _GEN_32 & _GEN_461;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1262 = _GEN_32 & _GEN_463;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1263 = _GEN_32 & _GEN_465;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1264 = _GEN_32 & _GEN_467;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1265 = _GEN_32 & _GEN_469;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1266 = _GEN_32 & _GEN_471;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1267 = _GEN_32 & _GEN_473;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1268 =
      _GEN_32 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1269 = _GEN_476 | _GEN_1237;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1270;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1271 = _GEN_479 | _GEN_1238;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1272;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1273 = _GEN_482 | _GEN_1239;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1274;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1275 = _GEN_485 | _GEN_1240;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1276;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1277 = _GEN_488 | _GEN_1241;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1278;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1279 = _GEN_491 | _GEN_1242;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1280;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1281 = _GEN_494 | _GEN_1243;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1282;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1283 = _GEN_497 | _GEN_1244;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1284;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1285 = _GEN_500 | _GEN_1245;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1286;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1287 = _GEN_503 | _GEN_1246;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1288;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1289 = _GEN_506 | _GEN_1247;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1290;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1291 = _GEN_509 | _GEN_1248;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1292;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1293 = _GEN_512 | _GEN_1249;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1294;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1295 = _GEN_515 | _GEN_1250;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1296;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1297 = _GEN_518 | _GEN_1251;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1298;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1299 = _GEN_521 | _GEN_1252;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1300;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1301 = _GEN_524 | _GEN_1253;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1302;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1303 = _GEN_527 | _GEN_1254;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1304;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1305 = _GEN_530 | _GEN_1255;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1306;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1307 = _GEN_533 | _GEN_1256;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1308;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1309 = _GEN_536 | _GEN_1257;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1310;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1311 = _GEN_539 | _GEN_1258;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1312;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1313 = _GEN_542 | _GEN_1259;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1314;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1315 = _GEN_545 | _GEN_1260;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1316;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1317 = _GEN_548 | _GEN_1261;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1318;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1319 = _GEN_551 | _GEN_1262;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1320;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1321 = _GEN_554 | _GEN_1263;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1322;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1323 = _GEN_557 | _GEN_1264;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1324;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1325 = _GEN_560 | _GEN_1265;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1326;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1327 = _GEN_563 | _GEN_1266;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1328;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1329 = _GEN_566 | _GEN_1267;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1330;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1331 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1268;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1332;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1333;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1334;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1335;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1336;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1337;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1338;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1339;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1340;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1341;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1342;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1343;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1344;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1345;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1346;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1347;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1348;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1349;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1350;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1351;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1352;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1353;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1354;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1355;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1356;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1357;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1358;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1359;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1360;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1361;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1362;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1363;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1364;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1365 = _GEN_34 & _GEN_603;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1366 = _GEN_34 & _GEN_605;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1367 = _GEN_34 & _GEN_607;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1368 = _GEN_34 & _GEN_609;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1369 = _GEN_34 & _GEN_611;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1370 = _GEN_34 & _GEN_613;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1371 = _GEN_34 & _GEN_615;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1372 = _GEN_34 & _GEN_617;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1373 = _GEN_34 & _GEN_619;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1374 = _GEN_34 & _GEN_621;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1375 = _GEN_34 & _GEN_623;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1376 = _GEN_34 & _GEN_625;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1377 = _GEN_34 & _GEN_627;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1378 = _GEN_34 & _GEN_629;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1379 = _GEN_34 & _GEN_631;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1380 = _GEN_34 & _GEN_633;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1381 = _GEN_34 & _GEN_635;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1382 = _GEN_34 & _GEN_637;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1383 = _GEN_34 & _GEN_639;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1384 = _GEN_34 & _GEN_641;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1385 = _GEN_34 & _GEN_643;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1386 = _GEN_34 & _GEN_645;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1387 = _GEN_34 & _GEN_647;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1388 = _GEN_34 & _GEN_649;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1389 = _GEN_34 & _GEN_651;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1390 = _GEN_34 & _GEN_653;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1391 = _GEN_34 & _GEN_655;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1392 = _GEN_34 & _GEN_657;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1393 = _GEN_34 & _GEN_659;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1394 = _GEN_34 & _GEN_661;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1395 = _GEN_34 & _GEN_663;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1396 =
      _GEN_34 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1397 = _GEN_666 | _GEN_1365;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1398;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1399 = _GEN_669 | _GEN_1366;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1400;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1401 = _GEN_672 | _GEN_1367;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1402;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1403 = _GEN_675 | _GEN_1368;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1404;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1405 = _GEN_678 | _GEN_1369;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1406;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1407 = _GEN_681 | _GEN_1370;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1408;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1409 = _GEN_684 | _GEN_1371;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1410;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1411 = _GEN_687 | _GEN_1372;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1412;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1413 = _GEN_690 | _GEN_1373;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1414;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1415 = _GEN_693 | _GEN_1374;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1416;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1417 = _GEN_696 | _GEN_1375;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1418;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1419 = _GEN_699 | _GEN_1376;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1420;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1421 = _GEN_702 | _GEN_1377;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1422;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1423 = _GEN_705 | _GEN_1378;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1424;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1425 = _GEN_708 | _GEN_1379;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1426;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1427 = _GEN_711 | _GEN_1380;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1428;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1429 = _GEN_714 | _GEN_1381;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1430;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1431 = _GEN_717 | _GEN_1382;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1432;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1433 = _GEN_720 | _GEN_1383;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1434;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1435 = _GEN_723 | _GEN_1384;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1436;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1437 = _GEN_726 | _GEN_1385;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1438;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1439 = _GEN_729 | _GEN_1386;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1440;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1441 = _GEN_732 | _GEN_1387;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1442;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1443 = _GEN_735 | _GEN_1388;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1444;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1445 = _GEN_738 | _GEN_1389;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1446;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1447 = _GEN_741 | _GEN_1390;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1448;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1449 = _GEN_744 | _GEN_1391;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1450;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1451 = _GEN_747 | _GEN_1392;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1452;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1453 = _GEN_750 | _GEN_1393;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1454;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1455 = _GEN_753 | _GEN_1394;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1456;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1457 = _GEN_756 | _GEN_1395;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1458;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1459 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1396;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1460;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1461;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1462;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1463;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1464;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1465;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1466;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1467;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1468;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1469;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1470;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1471;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1472;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1473;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1474;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1475;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1476;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1477;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1478;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1479;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1480;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1481;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1482;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1483;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1484;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1485;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1486;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1487;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1488;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1489;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1490;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1491;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1492;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1493;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1494;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1495;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1496;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1497;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1498;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1499;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1500;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1501;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1502;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1503;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1504;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1505;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1506;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1507;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1508;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1509;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1510;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1511;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1512;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1513;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1514;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1515;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1516;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1517;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1518;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1519;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1520;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1521;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1522;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1523;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1524;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_1525;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1526;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1527;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1528;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1529;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1530;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1531;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1532;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1533;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1534;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1535;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1536;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1537;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1538;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1539;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1540;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1541;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1542;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1543;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1544;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1545;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1546;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1547;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1548;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1549;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1550;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1551;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1552;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1553;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1554;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1555;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_1556;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [15:0]      _GEN_1557;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1558;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1559;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1560;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1561;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1562;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1563;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1564;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1565;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1566;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1567;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1568;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1569;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1570;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1571;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1572;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1573;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1574;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1575;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1576;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1577;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1578;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1579;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1580;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1581;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1582;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1583;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1584;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1585;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1586;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1587;	// util.scala:118:51
    automatic logic [15:0]      _GEN_1588;	// util.scala:118:51
    automatic logic             _GEN_1589;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1590;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1591;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1592;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1593;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1594;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1595;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1596;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1597;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1598;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1599;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1600;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1601;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1602;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1603;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1604;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1605;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1606;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1607;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1608;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1609;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1610;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1611;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1612;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1613;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1614;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1615;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1616;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1617;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1618;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1619;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _GEN_1620;	// rob.scala:307:32, :323:29, :324:31
    automatic logic             _rob_bsy_T_4 =
      io_enq_uops_2_is_fence | io_enq_uops_2_is_fencei;	// rob.scala:325:60
    automatic logic             _GEN_1621;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1622;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1623;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1624;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1625;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1626;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1627;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1628;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1629;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1630;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1631;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1632;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1633;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1634;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1635;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1636;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1637;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1638;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1639;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1640;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1641;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1642;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1643;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1644;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1645;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1646;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1647;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1648;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1649;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1650;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1651;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _GEN_1652;	// rob.scala:308:28, :323:29, :325:31
    automatic logic             _rob_unsafe_T_14 =
      io_enq_uops_2_uses_ldq | io_enq_uops_2_uses_stq & ~io_enq_uops_2_is_fence
      | io_enq_uops_2_is_br | io_enq_uops_2_is_jalr;	// micro-op.scala:152:{48,51,71}
    automatic logic             _GEN_1653;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1654;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1655;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1656;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1657;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1658;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1659;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1660;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1661;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1662;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1663;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1664;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1665;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1666;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1667;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1668;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1669;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1670;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1671;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1672;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1673;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1674;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1675;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1676;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1677;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1678;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1679;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1680;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1681;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1682;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1683;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1684;	// rob.scala:309:28, :323:29, :327:31
    automatic logic             _GEN_1685 = _GEN_60 & _GEN_223;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1686 = _GEN_60 & _GEN_225;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1687 = _GEN_60 & _GEN_227;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1688 = _GEN_60 & _GEN_229;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1689 = _GEN_60 & _GEN_231;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1690 = _GEN_60 & _GEN_233;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1691 = _GEN_60 & _GEN_235;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1692 = _GEN_60 & _GEN_237;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1693 = _GEN_60 & _GEN_239;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1694 = _GEN_60 & _GEN_241;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1695 = _GEN_60 & _GEN_243;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1696 = _GEN_60 & _GEN_245;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1697 = _GEN_60 & _GEN_247;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1698 = _GEN_60 & _GEN_249;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1699 = _GEN_60 & _GEN_251;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1700 = _GEN_60 & _GEN_253;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1701 = _GEN_60 & _GEN_255;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1702 = _GEN_60 & _GEN_257;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1703 = _GEN_60 & _GEN_259;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1704 = _GEN_60 & _GEN_261;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1705 = _GEN_60 & _GEN_263;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1706 = _GEN_60 & _GEN_265;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1707 = _GEN_60 & _GEN_267;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1708 = _GEN_60 & _GEN_269;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1709 = _GEN_60 & _GEN_271;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1710 = _GEN_60 & _GEN_273;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1711 = _GEN_60 & _GEN_275;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1712 = _GEN_60 & _GEN_277;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1713 = _GEN_60 & _GEN_279;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1714 = _GEN_60 & _GEN_281;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1715 = _GEN_60 & _GEN_283;	// rob.scala:323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1716 =
      _GEN_60 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :323:29, :346:{27,69}, :347:31
    automatic logic             _GEN_1717 = _GEN_286 | _GEN_1685;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1718;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1719 = _GEN_289 | _GEN_1686;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1720;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1721 = _GEN_292 | _GEN_1687;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1722;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1723 = _GEN_295 | _GEN_1688;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1724;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1725 = _GEN_298 | _GEN_1689;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1726;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1727 = _GEN_301 | _GEN_1690;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1728;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1729 = _GEN_304 | _GEN_1691;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1730;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1731 = _GEN_307 | _GEN_1692;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1732;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1733 = _GEN_310 | _GEN_1693;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1734;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1735 = _GEN_313 | _GEN_1694;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1736;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1737 = _GEN_316 | _GEN_1695;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1738;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1739 = _GEN_319 | _GEN_1696;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1740;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1741 = _GEN_322 | _GEN_1697;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1742;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1743 = _GEN_325 | _GEN_1698;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1744;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1745 = _GEN_328 | _GEN_1699;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1746;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1747 = _GEN_331 | _GEN_1700;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1748;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1749 = _GEN_334 | _GEN_1701;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1750;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1751 = _GEN_337 | _GEN_1702;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1752;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1753 = _GEN_340 | _GEN_1703;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1754;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1755 = _GEN_343 | _GEN_1704;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1756;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1757 = _GEN_346 | _GEN_1705;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1758;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1759 = _GEN_349 | _GEN_1706;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1760;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1761 = _GEN_352 | _GEN_1707;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1762;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1763 = _GEN_355 | _GEN_1708;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1764;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1765 = _GEN_358 | _GEN_1709;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1766;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1767 = _GEN_361 | _GEN_1710;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1768;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1769 = _GEN_364 | _GEN_1711;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1770;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1771 = _GEN_367 | _GEN_1712;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1772;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1773 = _GEN_370 | _GEN_1713;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1774;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1775 = _GEN_373 | _GEN_1714;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1776;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1777 = _GEN_376 | _GEN_1715;	// rob.scala:323:29, :346:69, :347:31
    automatic logic             _GEN_1778;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1779 =
      (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_1716;	// rob.scala:236:31, :268:25, :323:29, :346:69, :347:31
    automatic logic             _GEN_1780;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1781;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1782;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1783;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1784;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1785;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1786;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1787;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1788;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1789;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1790;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1791;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1792;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1793;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1794;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1795;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1796;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1797;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1798;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1799;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1800;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1801;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1802;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1803;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1804;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1805;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1806;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1807;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1808;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1809;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1810;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1811;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1812;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1813 = _GEN_62 & _GEN_413;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1814 = _GEN_62 & _GEN_415;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1815 = _GEN_62 & _GEN_417;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1816 = _GEN_62 & _GEN_419;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1817 = _GEN_62 & _GEN_421;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1818 = _GEN_62 & _GEN_423;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1819 = _GEN_62 & _GEN_425;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1820 = _GEN_62 & _GEN_427;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1821 = _GEN_62 & _GEN_429;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1822 = _GEN_62 & _GEN_431;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1823 = _GEN_62 & _GEN_433;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1824 = _GEN_62 & _GEN_435;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1825 = _GEN_62 & _GEN_437;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1826 = _GEN_62 & _GEN_439;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1827 = _GEN_62 & _GEN_441;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1828 = _GEN_62 & _GEN_443;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1829 = _GEN_62 & _GEN_445;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1830 = _GEN_62 & _GEN_447;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1831 = _GEN_62 & _GEN_449;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1832 = _GEN_62 & _GEN_451;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1833 = _GEN_62 & _GEN_453;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1834 = _GEN_62 & _GEN_455;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1835 = _GEN_62 & _GEN_457;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1836 = _GEN_62 & _GEN_459;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1837 = _GEN_62 & _GEN_461;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1838 = _GEN_62 & _GEN_463;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1839 = _GEN_62 & _GEN_465;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1840 = _GEN_62 & _GEN_467;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1841 = _GEN_62 & _GEN_469;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1842 = _GEN_62 & _GEN_471;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1843 = _GEN_62 & _GEN_473;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1844 =
      _GEN_62 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1845 = _GEN_476 | _GEN_1813;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1846;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1847 = _GEN_479 | _GEN_1814;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1848;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1849 = _GEN_482 | _GEN_1815;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1850;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1851 = _GEN_485 | _GEN_1816;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1852;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1853 = _GEN_488 | _GEN_1817;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1854;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1855 = _GEN_491 | _GEN_1818;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1856;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1857 = _GEN_494 | _GEN_1819;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1858;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1859 = _GEN_497 | _GEN_1820;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1860;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1861 = _GEN_500 | _GEN_1821;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1862;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1863 = _GEN_503 | _GEN_1822;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1864;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1865 = _GEN_506 | _GEN_1823;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1866;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1867 = _GEN_509 | _GEN_1824;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1868;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1869 = _GEN_512 | _GEN_1825;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1870;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1871 = _GEN_515 | _GEN_1826;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1872;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1873 = _GEN_518 | _GEN_1827;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1874;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1875 = _GEN_521 | _GEN_1828;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1876;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1877 = _GEN_524 | _GEN_1829;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1878;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1879 = _GEN_527 | _GEN_1830;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1880;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1881 = _GEN_530 | _GEN_1831;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1882;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1883 = _GEN_533 | _GEN_1832;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1884;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1885 = _GEN_536 | _GEN_1833;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1886;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1887 = _GEN_539 | _GEN_1834;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1888;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1889 = _GEN_542 | _GEN_1835;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1890;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1891 = _GEN_545 | _GEN_1836;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1892;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1893 = _GEN_548 | _GEN_1837;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1894;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1895 = _GEN_551 | _GEN_1838;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1896;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1897 = _GEN_554 | _GEN_1839;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1898;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1899 = _GEN_557 | _GEN_1840;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1900;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1901 = _GEN_560 | _GEN_1841;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1902;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1903 = _GEN_563 | _GEN_1842;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1904;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1905 = _GEN_566 | _GEN_1843;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1906;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1907 =
      (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1844;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_1908;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1909;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1910;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1911;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1912;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1913;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1914;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1915;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1916;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1917;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1918;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1919;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1920;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1921;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1922;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1923;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1924;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1925;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1926;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1927;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1928;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1929;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1930;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1931;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1932;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1933;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1934;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1935;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1936;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1937;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1938;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1939;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1940;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_1941 = _GEN_64 & _GEN_603;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1942 = _GEN_64 & _GEN_605;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1943 = _GEN_64 & _GEN_607;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1944 = _GEN_64 & _GEN_609;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1945 = _GEN_64 & _GEN_611;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1946 = _GEN_64 & _GEN_613;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1947 = _GEN_64 & _GEN_615;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1948 = _GEN_64 & _GEN_617;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1949 = _GEN_64 & _GEN_619;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1950 = _GEN_64 & _GEN_621;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1951 = _GEN_64 & _GEN_623;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1952 = _GEN_64 & _GEN_625;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1953 = _GEN_64 & _GEN_627;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1954 = _GEN_64 & _GEN_629;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1955 = _GEN_64 & _GEN_631;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1956 = _GEN_64 & _GEN_633;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1957 = _GEN_64 & _GEN_635;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1958 = _GEN_64 & _GEN_637;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1959 = _GEN_64 & _GEN_639;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1960 = _GEN_64 & _GEN_641;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1961 = _GEN_64 & _GEN_643;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1962 = _GEN_64 & _GEN_645;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1963 = _GEN_64 & _GEN_647;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1964 = _GEN_64 & _GEN_649;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1965 = _GEN_64 & _GEN_651;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1966 = _GEN_64 & _GEN_653;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1967 = _GEN_64 & _GEN_655;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1968 = _GEN_64 & _GEN_657;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1969 = _GEN_64 & _GEN_659;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1970 = _GEN_64 & _GEN_661;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1971 = _GEN_64 & _GEN_663;	// rob.scala:346:{27,69}, :347:31
    automatic logic             _GEN_1972 =
      _GEN_64 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));	// rob.scala:236:31, :268:25, :346:{27,69}, :347:31
    automatic logic             _GEN_1973 = _GEN_666 | _GEN_1941;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1974;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1975 = _GEN_669 | _GEN_1942;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1976;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1977 = _GEN_672 | _GEN_1943;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1978;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1979 = _GEN_675 | _GEN_1944;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1980;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1981 = _GEN_678 | _GEN_1945;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1982;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1983 = _GEN_681 | _GEN_1946;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1984;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1985 = _GEN_684 | _GEN_1947;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1986;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1987 = _GEN_687 | _GEN_1948;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1988;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1989 = _GEN_690 | _GEN_1949;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1990;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1991 = _GEN_693 | _GEN_1950;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1992;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1993 = _GEN_696 | _GEN_1951;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1994;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1995 = _GEN_699 | _GEN_1952;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1996;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1997 = _GEN_702 | _GEN_1953;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1998;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_1999 = _GEN_705 | _GEN_1954;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2000;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2001 = _GEN_708 | _GEN_1955;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2002;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2003 = _GEN_711 | _GEN_1956;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2004;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2005 = _GEN_714 | _GEN_1957;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2006;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2007 = _GEN_717 | _GEN_1958;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2008;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2009 = _GEN_720 | _GEN_1959;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2010;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2011 = _GEN_723 | _GEN_1960;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2012;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2013 = _GEN_726 | _GEN_1961;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2014;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2015 = _GEN_729 | _GEN_1962;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2016;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2017 = _GEN_732 | _GEN_1963;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2018;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2019 = _GEN_735 | _GEN_1964;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2020;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2021 = _GEN_738 | _GEN_1965;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2022;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2023 = _GEN_741 | _GEN_1966;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2024;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2025 = _GEN_744 | _GEN_1967;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2026;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2027 = _GEN_747 | _GEN_1968;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2028;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2029 = _GEN_750 | _GEN_1969;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2030;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2031 = _GEN_753 | _GEN_1970;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2032;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2033 = _GEN_756 | _GEN_1971;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2034;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2035 =
      (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1972;	// rob.scala:236:31, :268:25, :346:69, :347:31
    automatic logic             _GEN_2036;	// rob.scala:346:69, :347:31
    automatic logic             _GEN_2037;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2038;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2039;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2040;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2041;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2042;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2043;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2044;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2045;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2046;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2047;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2048;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2049;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2050;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2051;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2052;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2053;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2054;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2055;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2056;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2057;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2058;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2059;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2060;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2061;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2062;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2063;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2064;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2065;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2066;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2067;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2068;	// rob.scala:346:69, :348:31
    automatic logic             _GEN_2069;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2070;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2071;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2072;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2073;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2074;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2075;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2076;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2077;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2078;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2079;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2080;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2081;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2082;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2083;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2084;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2085;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2086;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2087;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2088;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2089;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2090;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2091;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2092;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2093;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2094;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2095;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2096;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2097;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2098;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2099;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2100;	// rob.scala:346:69, :361:75, :363:26
    automatic logic             _GEN_2101;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2102;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2103;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2104;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2105;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2106;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2107;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2108;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2109;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2110;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2111;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2112;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2113;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2114;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2115;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2116;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2117;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2118;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2119;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2120;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2121;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2122;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2123;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2124;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2125;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2126;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2127;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2128;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2129;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2130;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2131;	// rob.scala:323:29, :433:20, :434:30
    automatic logic             _GEN_2132;	// rob.scala:323:29, :433:20, :434:30
    automatic logic [15:0]      _GEN_2133;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2134;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2135;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2136;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2137;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2138;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2139;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2140;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2141;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2142;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2143;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2144;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2145;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2146;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2147;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2148;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2149;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2150;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2151;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2152;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2153;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2154;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2155;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2156;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2157;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2158;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2159;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2160;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2161;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2162;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2163;	// util.scala:118:51
    automatic logic [15:0]      _GEN_2164;	// util.scala:118:51
    automatic logic             enq_xcpts_0 = io_enq_valids_0 & io_enq_uops_0_exception;	// rob.scala:628:38
    automatic logic             enq_xcpts_1 = io_enq_valids_1 & io_enq_uops_1_exception;	// rob.scala:628:38
    automatic logic             _GEN_2165;	// rob.scala:631:47
    automatic logic             _GEN_2166;	// rob.scala:635:25
    automatic logic             _GEN_2167;	// rob.scala:641:30
    automatic logic [1:0]       idx;	// rob.scala:642:37
    automatic logic [3:0][15:0] _GEN_2168 =
      {{io_enq_uops_0_br_mask},
       {io_enq_uops_2_br_mask},
       {io_enq_uops_1_br_mask},
       {io_enq_uops_0_br_mask}};	// rob.scala:646:23
    automatic logic [15:0]      next_xcpt_uop_br_mask;	// rob.scala:625:17, :631:76, :632:27
    automatic logic [3:0]       _GEN_2169;	// rob.scala:865:98
    _GEN_96 = rob_tail == 5'h0;	// rob.scala:224:29, :228:29, :324:31
    _GEN_97 = io_enq_valids_0 & _GEN_96;	// rob.scala:307:32, :323:29, :324:31
    _GEN_98 = rob_tail == 5'h1;	// rob.scala:228:29, :324:31
    _GEN_99 = io_enq_valids_0 & _GEN_98;	// rob.scala:307:32, :323:29, :324:31
    _GEN_100 = rob_tail == 5'h2;	// rob.scala:228:29, :324:31
    _GEN_101 = io_enq_valids_0 & _GEN_100;	// rob.scala:307:32, :323:29, :324:31
    _GEN_102 = rob_tail == 5'h3;	// rob.scala:228:29, :324:31
    _GEN_103 = io_enq_valids_0 & _GEN_102;	// rob.scala:307:32, :323:29, :324:31
    _GEN_104 = rob_tail == 5'h4;	// rob.scala:228:29, :324:31
    _GEN_105 = io_enq_valids_0 & _GEN_104;	// rob.scala:307:32, :323:29, :324:31
    _GEN_106 = rob_tail == 5'h5;	// rob.scala:228:29, :324:31
    _GEN_107 = io_enq_valids_0 & _GEN_106;	// rob.scala:307:32, :323:29, :324:31
    _GEN_108 = rob_tail == 5'h6;	// rob.scala:228:29, :324:31
    _GEN_109 = io_enq_valids_0 & _GEN_108;	// rob.scala:307:32, :323:29, :324:31
    _GEN_110 = rob_tail == 5'h7;	// rob.scala:228:29, :324:31
    _GEN_111 = io_enq_valids_0 & _GEN_110;	// rob.scala:307:32, :323:29, :324:31
    _GEN_112 = rob_tail == 5'h8;	// rob.scala:228:29, :324:31
    _GEN_113 = io_enq_valids_0 & _GEN_112;	// rob.scala:307:32, :323:29, :324:31
    _GEN_114 = rob_tail == 5'h9;	// rob.scala:228:29, :324:31
    _GEN_115 = io_enq_valids_0 & _GEN_114;	// rob.scala:307:32, :323:29, :324:31
    _GEN_116 = rob_tail == 5'hA;	// rob.scala:228:29, :324:31
    _GEN_117 = io_enq_valids_0 & _GEN_116;	// rob.scala:307:32, :323:29, :324:31
    _GEN_118 = rob_tail == 5'hB;	// rob.scala:228:29, :324:31
    _GEN_119 = io_enq_valids_0 & _GEN_118;	// rob.scala:307:32, :323:29, :324:31
    _GEN_120 = rob_tail == 5'hC;	// rob.scala:228:29, :324:31
    _GEN_121 = io_enq_valids_0 & _GEN_120;	// rob.scala:307:32, :323:29, :324:31
    _GEN_122 = rob_tail == 5'hD;	// rob.scala:228:29, :324:31
    _GEN_123 = io_enq_valids_0 & _GEN_122;	// rob.scala:307:32, :323:29, :324:31
    _GEN_124 = rob_tail == 5'hE;	// rob.scala:228:29, :324:31
    _GEN_125 = io_enq_valids_0 & _GEN_124;	// rob.scala:307:32, :323:29, :324:31
    _GEN_126 = rob_tail == 5'hF;	// rob.scala:228:29, :324:31
    _GEN_127 = io_enq_valids_0 & _GEN_126;	// rob.scala:307:32, :323:29, :324:31
    _GEN_128 = rob_tail == 5'h10;	// rob.scala:228:29, :324:31
    _GEN_129 = io_enq_valids_0 & _GEN_128;	// rob.scala:307:32, :323:29, :324:31
    _GEN_130 = rob_tail == 5'h11;	// rob.scala:228:29, :324:31
    _GEN_131 = io_enq_valids_0 & _GEN_130;	// rob.scala:307:32, :323:29, :324:31
    _GEN_132 = rob_tail == 5'h12;	// rob.scala:228:29, :324:31
    _GEN_133 = io_enq_valids_0 & _GEN_132;	// rob.scala:307:32, :323:29, :324:31
    _GEN_134 = rob_tail == 5'h13;	// rob.scala:228:29, :324:31
    _GEN_135 = io_enq_valids_0 & _GEN_134;	// rob.scala:307:32, :323:29, :324:31
    _GEN_136 = rob_tail == 5'h14;	// rob.scala:228:29, :324:31
    _GEN_137 = io_enq_valids_0 & _GEN_136;	// rob.scala:307:32, :323:29, :324:31
    _GEN_138 = rob_tail == 5'h15;	// rob.scala:228:29, :324:31
    _GEN_139 = io_enq_valids_0 & _GEN_138;	// rob.scala:307:32, :323:29, :324:31
    _GEN_140 = rob_tail == 5'h16;	// rob.scala:228:29, :324:31
    _GEN_141 = io_enq_valids_0 & _GEN_140;	// rob.scala:307:32, :323:29, :324:31
    _GEN_142 = rob_tail == 5'h17;	// rob.scala:228:29, :324:31
    _GEN_143 = io_enq_valids_0 & _GEN_142;	// rob.scala:307:32, :323:29, :324:31
    _GEN_144 = rob_tail == 5'h18;	// rob.scala:228:29, :324:31
    _GEN_145 = io_enq_valids_0 & _GEN_144;	// rob.scala:307:32, :323:29, :324:31
    _GEN_146 = rob_tail == 5'h19;	// rob.scala:228:29, :324:31
    _GEN_147 = io_enq_valids_0 & _GEN_146;	// rob.scala:307:32, :323:29, :324:31
    _GEN_148 = rob_tail == 5'h1A;	// rob.scala:228:29, :324:31
    _GEN_149 = io_enq_valids_0 & _GEN_148;	// rob.scala:307:32, :323:29, :324:31
    _GEN_150 = rob_tail == 5'h1B;	// rob.scala:228:29, :324:31
    _GEN_151 = io_enq_valids_0 & _GEN_150;	// rob.scala:307:32, :323:29, :324:31
    _GEN_152 = rob_tail == 5'h1C;	// rob.scala:228:29, :324:31
    _GEN_153 = io_enq_valids_0 & _GEN_152;	// rob.scala:307:32, :323:29, :324:31
    _GEN_154 = rob_tail == 5'h1D;	// rob.scala:228:29, :324:31
    _GEN_155 = io_enq_valids_0 & _GEN_154;	// rob.scala:307:32, :323:29, :324:31
    _GEN_156 = rob_tail == 5'h1E;	// rob.scala:228:29, :324:31
    _GEN_157 = io_enq_valids_0 & _GEN_156;	// rob.scala:307:32, :323:29, :324:31
    _GEN_158 = io_enq_valids_0 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_159 = _GEN_97 ? ~_rob_bsy_T : rob_bsy_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_160 = _GEN_99 ? ~_rob_bsy_T : rob_bsy_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_161 = _GEN_101 ? ~_rob_bsy_T : rob_bsy_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_162 = _GEN_103 ? ~_rob_bsy_T : rob_bsy_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_163 = _GEN_105 ? ~_rob_bsy_T : rob_bsy_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_164 = _GEN_107 ? ~_rob_bsy_T : rob_bsy_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_165 = _GEN_109 ? ~_rob_bsy_T : rob_bsy_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_166 = _GEN_111 ? ~_rob_bsy_T : rob_bsy_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_167 = _GEN_113 ? ~_rob_bsy_T : rob_bsy_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_168 = _GEN_115 ? ~_rob_bsy_T : rob_bsy_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_169 = _GEN_117 ? ~_rob_bsy_T : rob_bsy_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_170 = _GEN_119 ? ~_rob_bsy_T : rob_bsy_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_171 = _GEN_121 ? ~_rob_bsy_T : rob_bsy_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_172 = _GEN_123 ? ~_rob_bsy_T : rob_bsy_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_173 = _GEN_125 ? ~_rob_bsy_T : rob_bsy_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_174 = _GEN_127 ? ~_rob_bsy_T : rob_bsy_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_175 = _GEN_129 ? ~_rob_bsy_T : rob_bsy_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_176 = _GEN_131 ? ~_rob_bsy_T : rob_bsy_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_177 = _GEN_133 ? ~_rob_bsy_T : rob_bsy_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_178 = _GEN_135 ? ~_rob_bsy_T : rob_bsy_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_179 = _GEN_137 ? ~_rob_bsy_T : rob_bsy_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_180 = _GEN_139 ? ~_rob_bsy_T : rob_bsy_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_181 = _GEN_141 ? ~_rob_bsy_T : rob_bsy_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_182 = _GEN_143 ? ~_rob_bsy_T : rob_bsy_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_183 = _GEN_145 ? ~_rob_bsy_T : rob_bsy_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_184 = _GEN_147 ? ~_rob_bsy_T : rob_bsy_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_185 = _GEN_149 ? ~_rob_bsy_T : rob_bsy_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_186 = _GEN_151 ? ~_rob_bsy_T : rob_bsy_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_187 = _GEN_153 ? ~_rob_bsy_T : rob_bsy_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_188 = _GEN_155 ? ~_rob_bsy_T : rob_bsy_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_189 = _GEN_157 ? ~_rob_bsy_T : rob_bsy_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_190 = _GEN_158 ? ~_rob_bsy_T : rob_bsy_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_191 = _GEN_97 ? _rob_unsafe_T_4 : rob_unsafe_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_192 = _GEN_99 ? _rob_unsafe_T_4 : rob_unsafe_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_193 = _GEN_101 ? _rob_unsafe_T_4 : rob_unsafe_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_194 = _GEN_103 ? _rob_unsafe_T_4 : rob_unsafe_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_195 = _GEN_105 ? _rob_unsafe_T_4 : rob_unsafe_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_196 = _GEN_107 ? _rob_unsafe_T_4 : rob_unsafe_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_197 = _GEN_109 ? _rob_unsafe_T_4 : rob_unsafe_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_198 = _GEN_111 ? _rob_unsafe_T_4 : rob_unsafe_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_199 = _GEN_113 ? _rob_unsafe_T_4 : rob_unsafe_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_200 = _GEN_115 ? _rob_unsafe_T_4 : rob_unsafe_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_201 = _GEN_117 ? _rob_unsafe_T_4 : rob_unsafe_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_202 = _GEN_119 ? _rob_unsafe_T_4 : rob_unsafe_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_203 = _GEN_121 ? _rob_unsafe_T_4 : rob_unsafe_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_204 = _GEN_123 ? _rob_unsafe_T_4 : rob_unsafe_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_205 = _GEN_125 ? _rob_unsafe_T_4 : rob_unsafe_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_206 = _GEN_127 ? _rob_unsafe_T_4 : rob_unsafe_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_207 = _GEN_129 ? _rob_unsafe_T_4 : rob_unsafe_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_208 = _GEN_131 ? _rob_unsafe_T_4 : rob_unsafe_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_209 = _GEN_133 ? _rob_unsafe_T_4 : rob_unsafe_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_210 = _GEN_135 ? _rob_unsafe_T_4 : rob_unsafe_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_211 = _GEN_137 ? _rob_unsafe_T_4 : rob_unsafe_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_212 = _GEN_139 ? _rob_unsafe_T_4 : rob_unsafe_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_213 = _GEN_141 ? _rob_unsafe_T_4 : rob_unsafe_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_214 = _GEN_143 ? _rob_unsafe_T_4 : rob_unsafe_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_215 = _GEN_145 ? _rob_unsafe_T_4 : rob_unsafe_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_216 = _GEN_147 ? _rob_unsafe_T_4 : rob_unsafe_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_217 = _GEN_149 ? _rob_unsafe_T_4 : rob_unsafe_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_218 = _GEN_151 ? _rob_unsafe_T_4 : rob_unsafe_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_219 = _GEN_153 ? _rob_unsafe_T_4 : rob_unsafe_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_220 = _GEN_155 ? _rob_unsafe_T_4 : rob_unsafe_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_221 = _GEN_157 ? _rob_unsafe_T_4 : rob_unsafe_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_222 = _GEN_158 ? _rob_unsafe_T_4 : rob_unsafe_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_288 = _GEN_1 ? ~_GEN_287 & _GEN_159 : ~_GEN_224 & _GEN_159;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_291 = _GEN_1 ? ~_GEN_290 & _GEN_160 : ~_GEN_226 & _GEN_160;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_294 = _GEN_1 ? ~_GEN_293 & _GEN_161 : ~_GEN_228 & _GEN_161;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_297 = _GEN_1 ? ~_GEN_296 & _GEN_162 : ~_GEN_230 & _GEN_162;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_300 = _GEN_1 ? ~_GEN_299 & _GEN_163 : ~_GEN_232 & _GEN_163;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_303 = _GEN_1 ? ~_GEN_302 & _GEN_164 : ~_GEN_234 & _GEN_164;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_306 = _GEN_1 ? ~_GEN_305 & _GEN_165 : ~_GEN_236 & _GEN_165;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_309 = _GEN_1 ? ~_GEN_308 & _GEN_166 : ~_GEN_238 & _GEN_166;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_312 = _GEN_1 ? ~_GEN_311 & _GEN_167 : ~_GEN_240 & _GEN_167;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_315 = _GEN_1 ? ~_GEN_314 & _GEN_168 : ~_GEN_242 & _GEN_168;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_318 = _GEN_1 ? ~_GEN_317 & _GEN_169 : ~_GEN_244 & _GEN_169;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_321 = _GEN_1 ? ~_GEN_320 & _GEN_170 : ~_GEN_246 & _GEN_170;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_324 = _GEN_1 ? ~_GEN_323 & _GEN_171 : ~_GEN_248 & _GEN_171;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_327 = _GEN_1 ? ~_GEN_326 & _GEN_172 : ~_GEN_250 & _GEN_172;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_330 = _GEN_1 ? ~_GEN_329 & _GEN_173 : ~_GEN_252 & _GEN_173;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_333 = _GEN_1 ? ~_GEN_332 & _GEN_174 : ~_GEN_254 & _GEN_174;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_336 = _GEN_1 ? ~_GEN_335 & _GEN_175 : ~_GEN_256 & _GEN_175;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_339 = _GEN_1 ? ~_GEN_338 & _GEN_176 : ~_GEN_258 & _GEN_176;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_342 = _GEN_1 ? ~_GEN_341 & _GEN_177 : ~_GEN_260 & _GEN_177;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_345 = _GEN_1 ? ~_GEN_344 & _GEN_178 : ~_GEN_262 & _GEN_178;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_348 = _GEN_1 ? ~_GEN_347 & _GEN_179 : ~_GEN_264 & _GEN_179;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_351 = _GEN_1 ? ~_GEN_350 & _GEN_180 : ~_GEN_266 & _GEN_180;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_354 = _GEN_1 ? ~_GEN_353 & _GEN_181 : ~_GEN_268 & _GEN_181;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_357 = _GEN_1 ? ~_GEN_356 & _GEN_182 : ~_GEN_270 & _GEN_182;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_360 = _GEN_1 ? ~_GEN_359 & _GEN_183 : ~_GEN_272 & _GEN_183;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_363 = _GEN_1 ? ~_GEN_362 & _GEN_184 : ~_GEN_274 & _GEN_184;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_366 = _GEN_1 ? ~_GEN_365 & _GEN_185 : ~_GEN_276 & _GEN_185;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_369 = _GEN_1 ? ~_GEN_368 & _GEN_186 : ~_GEN_278 & _GEN_186;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_372 = _GEN_1 ? ~_GEN_371 & _GEN_187 : ~_GEN_280 & _GEN_187;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_375 = _GEN_1 ? ~_GEN_374 & _GEN_188 : ~_GEN_282 & _GEN_188;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_378 = _GEN_1 ? ~_GEN_377 & _GEN_189 : ~_GEN_284 & _GEN_189;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_380 = _GEN_1 ? ~_GEN_379 & _GEN_190 : ~_GEN_285 & _GEN_190;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_381 = _GEN_1 ? ~_GEN_287 & _GEN_191 : ~_GEN_224 & _GEN_191;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_382 = _GEN_1 ? ~_GEN_290 & _GEN_192 : ~_GEN_226 & _GEN_192;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_383 = _GEN_1 ? ~_GEN_293 & _GEN_193 : ~_GEN_228 & _GEN_193;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_384 = _GEN_1 ? ~_GEN_296 & _GEN_194 : ~_GEN_230 & _GEN_194;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_385 = _GEN_1 ? ~_GEN_299 & _GEN_195 : ~_GEN_232 & _GEN_195;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_386 = _GEN_1 ? ~_GEN_302 & _GEN_196 : ~_GEN_234 & _GEN_196;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_387 = _GEN_1 ? ~_GEN_305 & _GEN_197 : ~_GEN_236 & _GEN_197;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_388 = _GEN_1 ? ~_GEN_308 & _GEN_198 : ~_GEN_238 & _GEN_198;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_389 = _GEN_1 ? ~_GEN_311 & _GEN_199 : ~_GEN_240 & _GEN_199;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_390 = _GEN_1 ? ~_GEN_314 & _GEN_200 : ~_GEN_242 & _GEN_200;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_391 = _GEN_1 ? ~_GEN_317 & _GEN_201 : ~_GEN_244 & _GEN_201;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_392 = _GEN_1 ? ~_GEN_320 & _GEN_202 : ~_GEN_246 & _GEN_202;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_393 = _GEN_1 ? ~_GEN_323 & _GEN_203 : ~_GEN_248 & _GEN_203;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_394 = _GEN_1 ? ~_GEN_326 & _GEN_204 : ~_GEN_250 & _GEN_204;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_395 = _GEN_1 ? ~_GEN_329 & _GEN_205 : ~_GEN_252 & _GEN_205;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_396 = _GEN_1 ? ~_GEN_332 & _GEN_206 : ~_GEN_254 & _GEN_206;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_397 = _GEN_1 ? ~_GEN_335 & _GEN_207 : ~_GEN_256 & _GEN_207;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_398 = _GEN_1 ? ~_GEN_338 & _GEN_208 : ~_GEN_258 & _GEN_208;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_399 = _GEN_1 ? ~_GEN_341 & _GEN_209 : ~_GEN_260 & _GEN_209;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_400 = _GEN_1 ? ~_GEN_344 & _GEN_210 : ~_GEN_262 & _GEN_210;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_401 = _GEN_1 ? ~_GEN_347 & _GEN_211 : ~_GEN_264 & _GEN_211;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_402 = _GEN_1 ? ~_GEN_350 & _GEN_212 : ~_GEN_266 & _GEN_212;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_403 = _GEN_1 ? ~_GEN_353 & _GEN_213 : ~_GEN_268 & _GEN_213;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_404 = _GEN_1 ? ~_GEN_356 & _GEN_214 : ~_GEN_270 & _GEN_214;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_405 = _GEN_1 ? ~_GEN_359 & _GEN_215 : ~_GEN_272 & _GEN_215;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_406 = _GEN_1 ? ~_GEN_362 & _GEN_216 : ~_GEN_274 & _GEN_216;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_407 = _GEN_1 ? ~_GEN_365 & _GEN_217 : ~_GEN_276 & _GEN_217;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_408 = _GEN_1 ? ~_GEN_368 & _GEN_218 : ~_GEN_278 & _GEN_218;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_409 = _GEN_1 ? ~_GEN_371 & _GEN_219 : ~_GEN_280 & _GEN_219;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_410 = _GEN_1 ? ~_GEN_374 & _GEN_220 : ~_GEN_282 & _GEN_220;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_411 = _GEN_1 ? ~_GEN_377 & _GEN_221 : ~_GEN_284 & _GEN_221;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_412 = _GEN_1 ? ~_GEN_379 & _GEN_222 : ~_GEN_285 & _GEN_222;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_478 = _GEN_3 ? ~_GEN_477 & _GEN_288 : ~_GEN_414 & _GEN_288;	// rob.scala:346:{27,69}, :347:31
    _GEN_481 = _GEN_3 ? ~_GEN_480 & _GEN_291 : ~_GEN_416 & _GEN_291;	// rob.scala:346:{27,69}, :347:31
    _GEN_484 = _GEN_3 ? ~_GEN_483 & _GEN_294 : ~_GEN_418 & _GEN_294;	// rob.scala:346:{27,69}, :347:31
    _GEN_487 = _GEN_3 ? ~_GEN_486 & _GEN_297 : ~_GEN_420 & _GEN_297;	// rob.scala:346:{27,69}, :347:31
    _GEN_490 = _GEN_3 ? ~_GEN_489 & _GEN_300 : ~_GEN_422 & _GEN_300;	// rob.scala:346:{27,69}, :347:31
    _GEN_493 = _GEN_3 ? ~_GEN_492 & _GEN_303 : ~_GEN_424 & _GEN_303;	// rob.scala:346:{27,69}, :347:31
    _GEN_496 = _GEN_3 ? ~_GEN_495 & _GEN_306 : ~_GEN_426 & _GEN_306;	// rob.scala:346:{27,69}, :347:31
    _GEN_499 = _GEN_3 ? ~_GEN_498 & _GEN_309 : ~_GEN_428 & _GEN_309;	// rob.scala:346:{27,69}, :347:31
    _GEN_502 = _GEN_3 ? ~_GEN_501 & _GEN_312 : ~_GEN_430 & _GEN_312;	// rob.scala:346:{27,69}, :347:31
    _GEN_505 = _GEN_3 ? ~_GEN_504 & _GEN_315 : ~_GEN_432 & _GEN_315;	// rob.scala:346:{27,69}, :347:31
    _GEN_508 = _GEN_3 ? ~_GEN_507 & _GEN_318 : ~_GEN_434 & _GEN_318;	// rob.scala:346:{27,69}, :347:31
    _GEN_511 = _GEN_3 ? ~_GEN_510 & _GEN_321 : ~_GEN_436 & _GEN_321;	// rob.scala:346:{27,69}, :347:31
    _GEN_514 = _GEN_3 ? ~_GEN_513 & _GEN_324 : ~_GEN_438 & _GEN_324;	// rob.scala:346:{27,69}, :347:31
    _GEN_517 = _GEN_3 ? ~_GEN_516 & _GEN_327 : ~_GEN_440 & _GEN_327;	// rob.scala:346:{27,69}, :347:31
    _GEN_520 = _GEN_3 ? ~_GEN_519 & _GEN_330 : ~_GEN_442 & _GEN_330;	// rob.scala:346:{27,69}, :347:31
    _GEN_523 = _GEN_3 ? ~_GEN_522 & _GEN_333 : ~_GEN_444 & _GEN_333;	// rob.scala:346:{27,69}, :347:31
    _GEN_526 = _GEN_3 ? ~_GEN_525 & _GEN_336 : ~_GEN_446 & _GEN_336;	// rob.scala:346:{27,69}, :347:31
    _GEN_529 = _GEN_3 ? ~_GEN_528 & _GEN_339 : ~_GEN_448 & _GEN_339;	// rob.scala:346:{27,69}, :347:31
    _GEN_532 = _GEN_3 ? ~_GEN_531 & _GEN_342 : ~_GEN_450 & _GEN_342;	// rob.scala:346:{27,69}, :347:31
    _GEN_535 = _GEN_3 ? ~_GEN_534 & _GEN_345 : ~_GEN_452 & _GEN_345;	// rob.scala:346:{27,69}, :347:31
    _GEN_538 = _GEN_3 ? ~_GEN_537 & _GEN_348 : ~_GEN_454 & _GEN_348;	// rob.scala:346:{27,69}, :347:31
    _GEN_541 = _GEN_3 ? ~_GEN_540 & _GEN_351 : ~_GEN_456 & _GEN_351;	// rob.scala:346:{27,69}, :347:31
    _GEN_544 = _GEN_3 ? ~_GEN_543 & _GEN_354 : ~_GEN_458 & _GEN_354;	// rob.scala:346:{27,69}, :347:31
    _GEN_547 = _GEN_3 ? ~_GEN_546 & _GEN_357 : ~_GEN_460 & _GEN_357;	// rob.scala:346:{27,69}, :347:31
    _GEN_550 = _GEN_3 ? ~_GEN_549 & _GEN_360 : ~_GEN_462 & _GEN_360;	// rob.scala:346:{27,69}, :347:31
    _GEN_553 = _GEN_3 ? ~_GEN_552 & _GEN_363 : ~_GEN_464 & _GEN_363;	// rob.scala:346:{27,69}, :347:31
    _GEN_556 = _GEN_3 ? ~_GEN_555 & _GEN_366 : ~_GEN_466 & _GEN_366;	// rob.scala:346:{27,69}, :347:31
    _GEN_559 = _GEN_3 ? ~_GEN_558 & _GEN_369 : ~_GEN_468 & _GEN_369;	// rob.scala:346:{27,69}, :347:31
    _GEN_562 = _GEN_3 ? ~_GEN_561 & _GEN_372 : ~_GEN_470 & _GEN_372;	// rob.scala:346:{27,69}, :347:31
    _GEN_565 = _GEN_3 ? ~_GEN_564 & _GEN_375 : ~_GEN_472 & _GEN_375;	// rob.scala:346:{27,69}, :347:31
    _GEN_568 = _GEN_3 ? ~_GEN_567 & _GEN_378 : ~_GEN_474 & _GEN_378;	// rob.scala:346:{27,69}, :347:31
    _GEN_570 = _GEN_3 ? ~_GEN_569 & _GEN_380 : ~_GEN_475 & _GEN_380;	// rob.scala:346:{27,69}, :347:31
    _GEN_571 = _GEN_3 ? ~_GEN_477 & _GEN_381 : ~_GEN_414 & _GEN_381;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_572 = _GEN_3 ? ~_GEN_480 & _GEN_382 : ~_GEN_416 & _GEN_382;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_573 = _GEN_3 ? ~_GEN_483 & _GEN_383 : ~_GEN_418 & _GEN_383;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_574 = _GEN_3 ? ~_GEN_486 & _GEN_384 : ~_GEN_420 & _GEN_384;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_575 = _GEN_3 ? ~_GEN_489 & _GEN_385 : ~_GEN_422 & _GEN_385;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_576 = _GEN_3 ? ~_GEN_492 & _GEN_386 : ~_GEN_424 & _GEN_386;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_577 = _GEN_3 ? ~_GEN_495 & _GEN_387 : ~_GEN_426 & _GEN_387;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_578 = _GEN_3 ? ~_GEN_498 & _GEN_388 : ~_GEN_428 & _GEN_388;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_579 = _GEN_3 ? ~_GEN_501 & _GEN_389 : ~_GEN_430 & _GEN_389;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_580 = _GEN_3 ? ~_GEN_504 & _GEN_390 : ~_GEN_432 & _GEN_390;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_581 = _GEN_3 ? ~_GEN_507 & _GEN_391 : ~_GEN_434 & _GEN_391;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_582 = _GEN_3 ? ~_GEN_510 & _GEN_392 : ~_GEN_436 & _GEN_392;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_583 = _GEN_3 ? ~_GEN_513 & _GEN_393 : ~_GEN_438 & _GEN_393;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_584 = _GEN_3 ? ~_GEN_516 & _GEN_394 : ~_GEN_440 & _GEN_394;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_585 = _GEN_3 ? ~_GEN_519 & _GEN_395 : ~_GEN_442 & _GEN_395;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_586 = _GEN_3 ? ~_GEN_522 & _GEN_396 : ~_GEN_444 & _GEN_396;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_587 = _GEN_3 ? ~_GEN_525 & _GEN_397 : ~_GEN_446 & _GEN_397;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_588 = _GEN_3 ? ~_GEN_528 & _GEN_398 : ~_GEN_448 & _GEN_398;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_589 = _GEN_3 ? ~_GEN_531 & _GEN_399 : ~_GEN_450 & _GEN_399;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_590 = _GEN_3 ? ~_GEN_534 & _GEN_400 : ~_GEN_452 & _GEN_400;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_591 = _GEN_3 ? ~_GEN_537 & _GEN_401 : ~_GEN_454 & _GEN_401;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_592 = _GEN_3 ? ~_GEN_540 & _GEN_402 : ~_GEN_456 & _GEN_402;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_593 = _GEN_3 ? ~_GEN_543 & _GEN_403 : ~_GEN_458 & _GEN_403;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_594 = _GEN_3 ? ~_GEN_546 & _GEN_404 : ~_GEN_460 & _GEN_404;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_595 = _GEN_3 ? ~_GEN_549 & _GEN_405 : ~_GEN_462 & _GEN_405;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_596 = _GEN_3 ? ~_GEN_552 & _GEN_406 : ~_GEN_464 & _GEN_406;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_597 = _GEN_3 ? ~_GEN_555 & _GEN_407 : ~_GEN_466 & _GEN_407;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_598 = _GEN_3 ? ~_GEN_558 & _GEN_408 : ~_GEN_468 & _GEN_408;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_599 = _GEN_3 ? ~_GEN_561 & _GEN_409 : ~_GEN_470 & _GEN_409;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_600 = _GEN_3 ? ~_GEN_564 & _GEN_410 : ~_GEN_472 & _GEN_410;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_601 = _GEN_3 ? ~_GEN_567 & _GEN_411 : ~_GEN_474 & _GEN_411;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_602 = _GEN_3 ? ~_GEN_569 & _GEN_412 : ~_GEN_475 & _GEN_412;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_668 = _GEN_5 ? ~_GEN_667 & _GEN_478 : ~_GEN_604 & _GEN_478;	// rob.scala:346:{27,69}, :347:31
    _GEN_671 = _GEN_5 ? ~_GEN_670 & _GEN_481 : ~_GEN_606 & _GEN_481;	// rob.scala:346:{27,69}, :347:31
    _GEN_674 = _GEN_5 ? ~_GEN_673 & _GEN_484 : ~_GEN_608 & _GEN_484;	// rob.scala:346:{27,69}, :347:31
    _GEN_677 = _GEN_5 ? ~_GEN_676 & _GEN_487 : ~_GEN_610 & _GEN_487;	// rob.scala:346:{27,69}, :347:31
    _GEN_680 = _GEN_5 ? ~_GEN_679 & _GEN_490 : ~_GEN_612 & _GEN_490;	// rob.scala:346:{27,69}, :347:31
    _GEN_683 = _GEN_5 ? ~_GEN_682 & _GEN_493 : ~_GEN_614 & _GEN_493;	// rob.scala:346:{27,69}, :347:31
    _GEN_686 = _GEN_5 ? ~_GEN_685 & _GEN_496 : ~_GEN_616 & _GEN_496;	// rob.scala:346:{27,69}, :347:31
    _GEN_689 = _GEN_5 ? ~_GEN_688 & _GEN_499 : ~_GEN_618 & _GEN_499;	// rob.scala:346:{27,69}, :347:31
    _GEN_692 = _GEN_5 ? ~_GEN_691 & _GEN_502 : ~_GEN_620 & _GEN_502;	// rob.scala:346:{27,69}, :347:31
    _GEN_695 = _GEN_5 ? ~_GEN_694 & _GEN_505 : ~_GEN_622 & _GEN_505;	// rob.scala:346:{27,69}, :347:31
    _GEN_698 = _GEN_5 ? ~_GEN_697 & _GEN_508 : ~_GEN_624 & _GEN_508;	// rob.scala:346:{27,69}, :347:31
    _GEN_701 = _GEN_5 ? ~_GEN_700 & _GEN_511 : ~_GEN_626 & _GEN_511;	// rob.scala:346:{27,69}, :347:31
    _GEN_704 = _GEN_5 ? ~_GEN_703 & _GEN_514 : ~_GEN_628 & _GEN_514;	// rob.scala:346:{27,69}, :347:31
    _GEN_707 = _GEN_5 ? ~_GEN_706 & _GEN_517 : ~_GEN_630 & _GEN_517;	// rob.scala:346:{27,69}, :347:31
    _GEN_710 = _GEN_5 ? ~_GEN_709 & _GEN_520 : ~_GEN_632 & _GEN_520;	// rob.scala:346:{27,69}, :347:31
    _GEN_713 = _GEN_5 ? ~_GEN_712 & _GEN_523 : ~_GEN_634 & _GEN_523;	// rob.scala:346:{27,69}, :347:31
    _GEN_716 = _GEN_5 ? ~_GEN_715 & _GEN_526 : ~_GEN_636 & _GEN_526;	// rob.scala:346:{27,69}, :347:31
    _GEN_719 = _GEN_5 ? ~_GEN_718 & _GEN_529 : ~_GEN_638 & _GEN_529;	// rob.scala:346:{27,69}, :347:31
    _GEN_722 = _GEN_5 ? ~_GEN_721 & _GEN_532 : ~_GEN_640 & _GEN_532;	// rob.scala:346:{27,69}, :347:31
    _GEN_725 = _GEN_5 ? ~_GEN_724 & _GEN_535 : ~_GEN_642 & _GEN_535;	// rob.scala:346:{27,69}, :347:31
    _GEN_728 = _GEN_5 ? ~_GEN_727 & _GEN_538 : ~_GEN_644 & _GEN_538;	// rob.scala:346:{27,69}, :347:31
    _GEN_731 = _GEN_5 ? ~_GEN_730 & _GEN_541 : ~_GEN_646 & _GEN_541;	// rob.scala:346:{27,69}, :347:31
    _GEN_734 = _GEN_5 ? ~_GEN_733 & _GEN_544 : ~_GEN_648 & _GEN_544;	// rob.scala:346:{27,69}, :347:31
    _GEN_737 = _GEN_5 ? ~_GEN_736 & _GEN_547 : ~_GEN_650 & _GEN_547;	// rob.scala:346:{27,69}, :347:31
    _GEN_740 = _GEN_5 ? ~_GEN_739 & _GEN_550 : ~_GEN_652 & _GEN_550;	// rob.scala:346:{27,69}, :347:31
    _GEN_743 = _GEN_5 ? ~_GEN_742 & _GEN_553 : ~_GEN_654 & _GEN_553;	// rob.scala:346:{27,69}, :347:31
    _GEN_746 = _GEN_5 ? ~_GEN_745 & _GEN_556 : ~_GEN_656 & _GEN_556;	// rob.scala:346:{27,69}, :347:31
    _GEN_749 = _GEN_5 ? ~_GEN_748 & _GEN_559 : ~_GEN_658 & _GEN_559;	// rob.scala:346:{27,69}, :347:31
    _GEN_752 = _GEN_5 ? ~_GEN_751 & _GEN_562 : ~_GEN_660 & _GEN_562;	// rob.scala:346:{27,69}, :347:31
    _GEN_755 = _GEN_5 ? ~_GEN_754 & _GEN_565 : ~_GEN_662 & _GEN_565;	// rob.scala:346:{27,69}, :347:31
    _GEN_758 = _GEN_5 ? ~_GEN_757 & _GEN_568 : ~_GEN_664 & _GEN_568;	// rob.scala:346:{27,69}, :347:31
    _GEN_760 = _GEN_5 ? ~_GEN_759 & _GEN_570 : ~_GEN_665 & _GEN_570;	// rob.scala:346:{27,69}, :347:31
    _GEN_761 = _GEN_5 ? ~_GEN_667 & _GEN_571 : ~_GEN_604 & _GEN_571;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_762 = _GEN_5 ? ~_GEN_670 & _GEN_572 : ~_GEN_606 & _GEN_572;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_763 = _GEN_5 ? ~_GEN_673 & _GEN_573 : ~_GEN_608 & _GEN_573;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_764 = _GEN_5 ? ~_GEN_676 & _GEN_574 : ~_GEN_610 & _GEN_574;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_765 = _GEN_5 ? ~_GEN_679 & _GEN_575 : ~_GEN_612 & _GEN_575;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_766 = _GEN_5 ? ~_GEN_682 & _GEN_576 : ~_GEN_614 & _GEN_576;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_767 = _GEN_5 ? ~_GEN_685 & _GEN_577 : ~_GEN_616 & _GEN_577;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_768 = _GEN_5 ? ~_GEN_688 & _GEN_578 : ~_GEN_618 & _GEN_578;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_769 = _GEN_5 ? ~_GEN_691 & _GEN_579 : ~_GEN_620 & _GEN_579;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_770 = _GEN_5 ? ~_GEN_694 & _GEN_580 : ~_GEN_622 & _GEN_580;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_771 = _GEN_5 ? ~_GEN_697 & _GEN_581 : ~_GEN_624 & _GEN_581;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_772 = _GEN_5 ? ~_GEN_700 & _GEN_582 : ~_GEN_626 & _GEN_582;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_773 = _GEN_5 ? ~_GEN_703 & _GEN_583 : ~_GEN_628 & _GEN_583;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_774 = _GEN_5 ? ~_GEN_706 & _GEN_584 : ~_GEN_630 & _GEN_584;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_775 = _GEN_5 ? ~_GEN_709 & _GEN_585 : ~_GEN_632 & _GEN_585;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_776 = _GEN_5 ? ~_GEN_712 & _GEN_586 : ~_GEN_634 & _GEN_586;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_777 = _GEN_5 ? ~_GEN_715 & _GEN_587 : ~_GEN_636 & _GEN_587;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_778 = _GEN_5 ? ~_GEN_718 & _GEN_588 : ~_GEN_638 & _GEN_588;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_779 = _GEN_5 ? ~_GEN_721 & _GEN_589 : ~_GEN_640 & _GEN_589;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_780 = _GEN_5 ? ~_GEN_724 & _GEN_590 : ~_GEN_642 & _GEN_590;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_781 = _GEN_5 ? ~_GEN_727 & _GEN_591 : ~_GEN_644 & _GEN_591;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_782 = _GEN_5 ? ~_GEN_730 & _GEN_592 : ~_GEN_646 & _GEN_592;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_783 = _GEN_5 ? ~_GEN_733 & _GEN_593 : ~_GEN_648 & _GEN_593;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_784 = _GEN_5 ? ~_GEN_736 & _GEN_594 : ~_GEN_650 & _GEN_594;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_785 = _GEN_5 ? ~_GEN_739 & _GEN_595 : ~_GEN_652 & _GEN_595;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_786 = _GEN_5 ? ~_GEN_742 & _GEN_596 : ~_GEN_654 & _GEN_596;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_787 = _GEN_5 ? ~_GEN_745 & _GEN_597 : ~_GEN_656 & _GEN_597;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_788 = _GEN_5 ? ~_GEN_748 & _GEN_598 : ~_GEN_658 & _GEN_598;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_789 = _GEN_5 ? ~_GEN_751 & _GEN_599 : ~_GEN_660 & _GEN_599;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_790 = _GEN_5 ? ~_GEN_754 & _GEN_600 : ~_GEN_662 & _GEN_600;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_791 = _GEN_5 ? ~_GEN_757 & _GEN_601 : ~_GEN_664 & _GEN_601;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_792 = _GEN_5 ? ~_GEN_759 & _GEN_602 : ~_GEN_665 & _GEN_602;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_794 = _GEN_6 & _GEN_793;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_796 = _GEN_6 & _GEN_795;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_798 = _GEN_6 & _GEN_797;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_800 = _GEN_6 & _GEN_799;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_802 = _GEN_6 & _GEN_801;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_804 = _GEN_6 & _GEN_803;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_806 = _GEN_6 & _GEN_805;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_808 = _GEN_6 & _GEN_807;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_810 = _GEN_6 & _GEN_809;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_812 = _GEN_6 & _GEN_811;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_814 = _GEN_6 & _GEN_813;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_816 = _GEN_6 & _GEN_815;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_818 = _GEN_6 & _GEN_817;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_820 = _GEN_6 & _GEN_819;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_822 = _GEN_6 & _GEN_821;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_824 = _GEN_6 & _GEN_823;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_826 = _GEN_6 & _GEN_825;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_828 = _GEN_6 & _GEN_827;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_830 = _GEN_6 & _GEN_829;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_832 = _GEN_6 & _GEN_831;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_834 = _GEN_6 & _GEN_833;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_836 = _GEN_6 & _GEN_835;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_838 = _GEN_6 & _GEN_837;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_840 = _GEN_6 & _GEN_839;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_842 = _GEN_6 & _GEN_841;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_844 = _GEN_6 & _GEN_843;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_846 = _GEN_6 & _GEN_845;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_848 = _GEN_6 & _GEN_847;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_850 = _GEN_6 & _GEN_849;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_852 = _GEN_6 & _GEN_851;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_854 = _GEN_6 & _GEN_853;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_855 = _GEN_6 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    _GEN_856 = io_lsu_clr_bsy_1_bits[6:2] == 5'h0;	// rob.scala:224:29, :236:31, :268:25, :363:26
    _GEN_857 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_858 = io_lsu_clr_bsy_1_bits[6:2] == 5'h2;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_859 = io_lsu_clr_bsy_1_bits[6:2] == 5'h3;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_860 = io_lsu_clr_bsy_1_bits[6:2] == 5'h4;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_861 = io_lsu_clr_bsy_1_bits[6:2] == 5'h5;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_862 = io_lsu_clr_bsy_1_bits[6:2] == 5'h6;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_863 = io_lsu_clr_bsy_1_bits[6:2] == 5'h7;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_864 = io_lsu_clr_bsy_1_bits[6:2] == 5'h8;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_865 = io_lsu_clr_bsy_1_bits[6:2] == 5'h9;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_866 = io_lsu_clr_bsy_1_bits[6:2] == 5'hA;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_867 = io_lsu_clr_bsy_1_bits[6:2] == 5'hB;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_868 = io_lsu_clr_bsy_1_bits[6:2] == 5'hC;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_869 = io_lsu_clr_bsy_1_bits[6:2] == 5'hD;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_870 = io_lsu_clr_bsy_1_bits[6:2] == 5'hE;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_871 = io_lsu_clr_bsy_1_bits[6:2] == 5'hF;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_872 = io_lsu_clr_bsy_1_bits[6:2] == 5'h10;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_873 = io_lsu_clr_bsy_1_bits[6:2] == 5'h11;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_874 = io_lsu_clr_bsy_1_bits[6:2] == 5'h12;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_875 = io_lsu_clr_bsy_1_bits[6:2] == 5'h13;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_876 = io_lsu_clr_bsy_1_bits[6:2] == 5'h14;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_877 = io_lsu_clr_bsy_1_bits[6:2] == 5'h15;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_878 = io_lsu_clr_bsy_1_bits[6:2] == 5'h16;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_879 = io_lsu_clr_bsy_1_bits[6:2] == 5'h17;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_880 = io_lsu_clr_bsy_1_bits[6:2] == 5'h18;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_881 = io_lsu_clr_bsy_1_bits[6:2] == 5'h19;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_882 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1A;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_883 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1B;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_884 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1C;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_885 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1D;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_886 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1E;	// rob.scala:236:31, :268:25, :324:31, :363:26
    _GEN_919 = rbk_row & _GEN_918;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_921 = rbk_row & _GEN_920;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_923 = rbk_row & _GEN_922;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_925 = rbk_row & _GEN_924;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_927 = rbk_row & _GEN_926;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_929 = rbk_row & _GEN_928;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_931 = rbk_row & _GEN_930;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_933 = rbk_row & _GEN_932;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_935 = rbk_row & _GEN_934;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_937 = rbk_row & _GEN_936;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_939 = rbk_row & _GEN_938;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_941 = rbk_row & _GEN_940;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_943 = rbk_row & _GEN_942;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_945 = rbk_row & _GEN_944;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_947 = rbk_row & _GEN_946;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_949 = rbk_row & _GEN_948;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_951 = rbk_row & _GEN_950;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_953 = rbk_row & _GEN_952;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_955 = rbk_row & _GEN_954;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_957 = rbk_row & _GEN_956;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_959 = rbk_row & _GEN_958;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_961 = rbk_row & _GEN_960;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_963 = rbk_row & _GEN_962;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_965 = rbk_row & _GEN_964;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_967 = rbk_row & _GEN_966;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_969 = rbk_row & _GEN_968;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_971 = rbk_row & _GEN_970;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_973 = rbk_row & _GEN_972;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_975 = rbk_row & _GEN_974;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_977 = rbk_row & _GEN_976;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_979 = rbk_row & _GEN_978;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_980 = rbk_row & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_981 = io_brupdate_b1_mispredict_mask & rob_uop_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_982 = io_brupdate_b1_mispredict_mask & rob_uop_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_983 = io_brupdate_b1_mispredict_mask & rob_uop_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_984 = io_brupdate_b1_mispredict_mask & rob_uop_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_985 = io_brupdate_b1_mispredict_mask & rob_uop_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_986 = io_brupdate_b1_mispredict_mask & rob_uop_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_987 = io_brupdate_b1_mispredict_mask & rob_uop_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_988 = io_brupdate_b1_mispredict_mask & rob_uop_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_989 = io_brupdate_b1_mispredict_mask & rob_uop_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_990 = io_brupdate_b1_mispredict_mask & rob_uop_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_991 = io_brupdate_b1_mispredict_mask & rob_uop_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_992 = io_brupdate_b1_mispredict_mask & rob_uop_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_993 = io_brupdate_b1_mispredict_mask & rob_uop_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_994 = io_brupdate_b1_mispredict_mask & rob_uop_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_995 = io_brupdate_b1_mispredict_mask & rob_uop_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_996 = io_brupdate_b1_mispredict_mask & rob_uop_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_997 = io_brupdate_b1_mispredict_mask & rob_uop_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_998 = io_brupdate_b1_mispredict_mask & rob_uop_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_999 = io_brupdate_b1_mispredict_mask & rob_uop_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1000 = io_brupdate_b1_mispredict_mask & rob_uop_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1001 = io_brupdate_b1_mispredict_mask & rob_uop_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1002 = io_brupdate_b1_mispredict_mask & rob_uop_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1003 = io_brupdate_b1_mispredict_mask & rob_uop_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1004 = io_brupdate_b1_mispredict_mask & rob_uop_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1005 = io_brupdate_b1_mispredict_mask & rob_uop_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1006 = io_brupdate_b1_mispredict_mask & rob_uop_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1007 = io_brupdate_b1_mispredict_mask & rob_uop_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1008 = io_brupdate_b1_mispredict_mask & rob_uop_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1009 = io_brupdate_b1_mispredict_mask & rob_uop_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1010 = io_brupdate_b1_mispredict_mask & rob_uop_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1011 = io_brupdate_b1_mispredict_mask & rob_uop_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1012 = io_brupdate_b1_mispredict_mask & rob_uop_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    rob_head_uses_ldq_0 = _GEN_21[rob_head];	// rob.scala:224:29, :411:25, :484:26
    _GEN_1013 = io_enq_valids_1 & _GEN_96;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1014 = io_enq_valids_1 & _GEN_98;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1015 = io_enq_valids_1 & _GEN_100;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1016 = io_enq_valids_1 & _GEN_102;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1017 = io_enq_valids_1 & _GEN_104;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1018 = io_enq_valids_1 & _GEN_106;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1019 = io_enq_valids_1 & _GEN_108;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1020 = io_enq_valids_1 & _GEN_110;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1021 = io_enq_valids_1 & _GEN_112;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1022 = io_enq_valids_1 & _GEN_114;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1023 = io_enq_valids_1 & _GEN_116;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1024 = io_enq_valids_1 & _GEN_118;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1025 = io_enq_valids_1 & _GEN_120;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1026 = io_enq_valids_1 & _GEN_122;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1027 = io_enq_valids_1 & _GEN_124;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1028 = io_enq_valids_1 & _GEN_126;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1029 = io_enq_valids_1 & _GEN_128;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1030 = io_enq_valids_1 & _GEN_130;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1031 = io_enq_valids_1 & _GEN_132;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1032 = io_enq_valids_1 & _GEN_134;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1033 = io_enq_valids_1 & _GEN_136;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1034 = io_enq_valids_1 & _GEN_138;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1035 = io_enq_valids_1 & _GEN_140;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1036 = io_enq_valids_1 & _GEN_142;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1037 = io_enq_valids_1 & _GEN_144;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1038 = io_enq_valids_1 & _GEN_146;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1039 = io_enq_valids_1 & _GEN_148;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1040 = io_enq_valids_1 & _GEN_150;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1041 = io_enq_valids_1 & _GEN_152;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1042 = io_enq_valids_1 & _GEN_154;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1043 = io_enq_valids_1 & _GEN_156;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1044 = io_enq_valids_1 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_1045 = _GEN_1013 ? ~_rob_bsy_T_2 : rob_bsy_1_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1046 = _GEN_1014 ? ~_rob_bsy_T_2 : rob_bsy_1_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1047 = _GEN_1015 ? ~_rob_bsy_T_2 : rob_bsy_1_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1048 = _GEN_1016 ? ~_rob_bsy_T_2 : rob_bsy_1_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1049 = _GEN_1017 ? ~_rob_bsy_T_2 : rob_bsy_1_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1050 = _GEN_1018 ? ~_rob_bsy_T_2 : rob_bsy_1_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1051 = _GEN_1019 ? ~_rob_bsy_T_2 : rob_bsy_1_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1052 = _GEN_1020 ? ~_rob_bsy_T_2 : rob_bsy_1_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1053 = _GEN_1021 ? ~_rob_bsy_T_2 : rob_bsy_1_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1054 = _GEN_1022 ? ~_rob_bsy_T_2 : rob_bsy_1_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1055 = _GEN_1023 ? ~_rob_bsy_T_2 : rob_bsy_1_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1056 = _GEN_1024 ? ~_rob_bsy_T_2 : rob_bsy_1_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1057 = _GEN_1025 ? ~_rob_bsy_T_2 : rob_bsy_1_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1058 = _GEN_1026 ? ~_rob_bsy_T_2 : rob_bsy_1_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1059 = _GEN_1027 ? ~_rob_bsy_T_2 : rob_bsy_1_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1060 = _GEN_1028 ? ~_rob_bsy_T_2 : rob_bsy_1_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1061 = _GEN_1029 ? ~_rob_bsy_T_2 : rob_bsy_1_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1062 = _GEN_1030 ? ~_rob_bsy_T_2 : rob_bsy_1_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1063 = _GEN_1031 ? ~_rob_bsy_T_2 : rob_bsy_1_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1064 = _GEN_1032 ? ~_rob_bsy_T_2 : rob_bsy_1_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1065 = _GEN_1033 ? ~_rob_bsy_T_2 : rob_bsy_1_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1066 = _GEN_1034 ? ~_rob_bsy_T_2 : rob_bsy_1_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1067 = _GEN_1035 ? ~_rob_bsy_T_2 : rob_bsy_1_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1068 = _GEN_1036 ? ~_rob_bsy_T_2 : rob_bsy_1_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1069 = _GEN_1037 ? ~_rob_bsy_T_2 : rob_bsy_1_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1070 = _GEN_1038 ? ~_rob_bsy_T_2 : rob_bsy_1_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1071 = _GEN_1039 ? ~_rob_bsy_T_2 : rob_bsy_1_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1072 = _GEN_1040 ? ~_rob_bsy_T_2 : rob_bsy_1_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1073 = _GEN_1041 ? ~_rob_bsy_T_2 : rob_bsy_1_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1074 = _GEN_1042 ? ~_rob_bsy_T_2 : rob_bsy_1_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1075 = _GEN_1043 ? ~_rob_bsy_T_2 : rob_bsy_1_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1076 = _GEN_1044 ? ~_rob_bsy_T_2 : rob_bsy_1_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1077 = _GEN_1013 ? _rob_unsafe_T_9 : rob_unsafe_1_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1078 = _GEN_1014 ? _rob_unsafe_T_9 : rob_unsafe_1_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1079 = _GEN_1015 ? _rob_unsafe_T_9 : rob_unsafe_1_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1080 = _GEN_1016 ? _rob_unsafe_T_9 : rob_unsafe_1_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1081 = _GEN_1017 ? _rob_unsafe_T_9 : rob_unsafe_1_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1082 = _GEN_1018 ? _rob_unsafe_T_9 : rob_unsafe_1_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1083 = _GEN_1019 ? _rob_unsafe_T_9 : rob_unsafe_1_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1084 = _GEN_1020 ? _rob_unsafe_T_9 : rob_unsafe_1_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1085 = _GEN_1021 ? _rob_unsafe_T_9 : rob_unsafe_1_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1086 = _GEN_1022 ? _rob_unsafe_T_9 : rob_unsafe_1_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1087 = _GEN_1023 ? _rob_unsafe_T_9 : rob_unsafe_1_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1088 = _GEN_1024 ? _rob_unsafe_T_9 : rob_unsafe_1_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1089 = _GEN_1025 ? _rob_unsafe_T_9 : rob_unsafe_1_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1090 = _GEN_1026 ? _rob_unsafe_T_9 : rob_unsafe_1_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1091 = _GEN_1027 ? _rob_unsafe_T_9 : rob_unsafe_1_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1092 = _GEN_1028 ? _rob_unsafe_T_9 : rob_unsafe_1_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1093 = _GEN_1029 ? _rob_unsafe_T_9 : rob_unsafe_1_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1094 = _GEN_1030 ? _rob_unsafe_T_9 : rob_unsafe_1_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1095 = _GEN_1031 ? _rob_unsafe_T_9 : rob_unsafe_1_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1096 = _GEN_1032 ? _rob_unsafe_T_9 : rob_unsafe_1_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1097 = _GEN_1033 ? _rob_unsafe_T_9 : rob_unsafe_1_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1098 = _GEN_1034 ? _rob_unsafe_T_9 : rob_unsafe_1_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1099 = _GEN_1035 ? _rob_unsafe_T_9 : rob_unsafe_1_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1100 = _GEN_1036 ? _rob_unsafe_T_9 : rob_unsafe_1_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1101 = _GEN_1037 ? _rob_unsafe_T_9 : rob_unsafe_1_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1102 = _GEN_1038 ? _rob_unsafe_T_9 : rob_unsafe_1_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1103 = _GEN_1039 ? _rob_unsafe_T_9 : rob_unsafe_1_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1104 = _GEN_1040 ? _rob_unsafe_T_9 : rob_unsafe_1_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1105 = _GEN_1041 ? _rob_unsafe_T_9 : rob_unsafe_1_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1106 = _GEN_1042 ? _rob_unsafe_T_9 : rob_unsafe_1_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1107 = _GEN_1043 ? _rob_unsafe_T_9 : rob_unsafe_1_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1108 = _GEN_1044 ? _rob_unsafe_T_9 : rob_unsafe_1_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1142 = _GEN_31 ? ~_GEN_1141 & _GEN_1045 : ~_GEN_1109 & _GEN_1045;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1144 = _GEN_31 ? ~_GEN_1143 & _GEN_1046 : ~_GEN_1110 & _GEN_1046;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1146 = _GEN_31 ? ~_GEN_1145 & _GEN_1047 : ~_GEN_1111 & _GEN_1047;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1148 = _GEN_31 ? ~_GEN_1147 & _GEN_1048 : ~_GEN_1112 & _GEN_1048;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1150 = _GEN_31 ? ~_GEN_1149 & _GEN_1049 : ~_GEN_1113 & _GEN_1049;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1152 = _GEN_31 ? ~_GEN_1151 & _GEN_1050 : ~_GEN_1114 & _GEN_1050;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1154 = _GEN_31 ? ~_GEN_1153 & _GEN_1051 : ~_GEN_1115 & _GEN_1051;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1156 = _GEN_31 ? ~_GEN_1155 & _GEN_1052 : ~_GEN_1116 & _GEN_1052;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1158 = _GEN_31 ? ~_GEN_1157 & _GEN_1053 : ~_GEN_1117 & _GEN_1053;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1160 = _GEN_31 ? ~_GEN_1159 & _GEN_1054 : ~_GEN_1118 & _GEN_1054;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1162 = _GEN_31 ? ~_GEN_1161 & _GEN_1055 : ~_GEN_1119 & _GEN_1055;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1164 = _GEN_31 ? ~_GEN_1163 & _GEN_1056 : ~_GEN_1120 & _GEN_1056;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1166 = _GEN_31 ? ~_GEN_1165 & _GEN_1057 : ~_GEN_1121 & _GEN_1057;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1168 = _GEN_31 ? ~_GEN_1167 & _GEN_1058 : ~_GEN_1122 & _GEN_1058;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1170 = _GEN_31 ? ~_GEN_1169 & _GEN_1059 : ~_GEN_1123 & _GEN_1059;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1172 = _GEN_31 ? ~_GEN_1171 & _GEN_1060 : ~_GEN_1124 & _GEN_1060;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1174 = _GEN_31 ? ~_GEN_1173 & _GEN_1061 : ~_GEN_1125 & _GEN_1061;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1176 = _GEN_31 ? ~_GEN_1175 & _GEN_1062 : ~_GEN_1126 & _GEN_1062;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1178 = _GEN_31 ? ~_GEN_1177 & _GEN_1063 : ~_GEN_1127 & _GEN_1063;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1180 = _GEN_31 ? ~_GEN_1179 & _GEN_1064 : ~_GEN_1128 & _GEN_1064;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1182 = _GEN_31 ? ~_GEN_1181 & _GEN_1065 : ~_GEN_1129 & _GEN_1065;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1184 = _GEN_31 ? ~_GEN_1183 & _GEN_1066 : ~_GEN_1130 & _GEN_1066;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1186 = _GEN_31 ? ~_GEN_1185 & _GEN_1067 : ~_GEN_1131 & _GEN_1067;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1188 = _GEN_31 ? ~_GEN_1187 & _GEN_1068 : ~_GEN_1132 & _GEN_1068;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1190 = _GEN_31 ? ~_GEN_1189 & _GEN_1069 : ~_GEN_1133 & _GEN_1069;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1192 = _GEN_31 ? ~_GEN_1191 & _GEN_1070 : ~_GEN_1134 & _GEN_1070;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1194 = _GEN_31 ? ~_GEN_1193 & _GEN_1071 : ~_GEN_1135 & _GEN_1071;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1196 = _GEN_31 ? ~_GEN_1195 & _GEN_1072 : ~_GEN_1136 & _GEN_1072;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1198 = _GEN_31 ? ~_GEN_1197 & _GEN_1073 : ~_GEN_1137 & _GEN_1073;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1200 = _GEN_31 ? ~_GEN_1199 & _GEN_1074 : ~_GEN_1138 & _GEN_1074;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1202 = _GEN_31 ? ~_GEN_1201 & _GEN_1075 : ~_GEN_1139 & _GEN_1075;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1204 = _GEN_31 ? ~_GEN_1203 & _GEN_1076 : ~_GEN_1140 & _GEN_1076;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1205 = _GEN_31 ? ~_GEN_1141 & _GEN_1077 : ~_GEN_1109 & _GEN_1077;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1206 = _GEN_31 ? ~_GEN_1143 & _GEN_1078 : ~_GEN_1110 & _GEN_1078;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1207 = _GEN_31 ? ~_GEN_1145 & _GEN_1079 : ~_GEN_1111 & _GEN_1079;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1208 = _GEN_31 ? ~_GEN_1147 & _GEN_1080 : ~_GEN_1112 & _GEN_1080;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1209 = _GEN_31 ? ~_GEN_1149 & _GEN_1081 : ~_GEN_1113 & _GEN_1081;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1210 = _GEN_31 ? ~_GEN_1151 & _GEN_1082 : ~_GEN_1114 & _GEN_1082;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1211 = _GEN_31 ? ~_GEN_1153 & _GEN_1083 : ~_GEN_1115 & _GEN_1083;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1212 = _GEN_31 ? ~_GEN_1155 & _GEN_1084 : ~_GEN_1116 & _GEN_1084;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1213 = _GEN_31 ? ~_GEN_1157 & _GEN_1085 : ~_GEN_1117 & _GEN_1085;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1214 = _GEN_31 ? ~_GEN_1159 & _GEN_1086 : ~_GEN_1118 & _GEN_1086;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1215 = _GEN_31 ? ~_GEN_1161 & _GEN_1087 : ~_GEN_1119 & _GEN_1087;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1216 = _GEN_31 ? ~_GEN_1163 & _GEN_1088 : ~_GEN_1120 & _GEN_1088;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1217 = _GEN_31 ? ~_GEN_1165 & _GEN_1089 : ~_GEN_1121 & _GEN_1089;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1218 = _GEN_31 ? ~_GEN_1167 & _GEN_1090 : ~_GEN_1122 & _GEN_1090;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1219 = _GEN_31 ? ~_GEN_1169 & _GEN_1091 : ~_GEN_1123 & _GEN_1091;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1220 = _GEN_31 ? ~_GEN_1171 & _GEN_1092 : ~_GEN_1124 & _GEN_1092;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1221 = _GEN_31 ? ~_GEN_1173 & _GEN_1093 : ~_GEN_1125 & _GEN_1093;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1222 = _GEN_31 ? ~_GEN_1175 & _GEN_1094 : ~_GEN_1126 & _GEN_1094;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1223 = _GEN_31 ? ~_GEN_1177 & _GEN_1095 : ~_GEN_1127 & _GEN_1095;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1224 = _GEN_31 ? ~_GEN_1179 & _GEN_1096 : ~_GEN_1128 & _GEN_1096;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1225 = _GEN_31 ? ~_GEN_1181 & _GEN_1097 : ~_GEN_1129 & _GEN_1097;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1226 = _GEN_31 ? ~_GEN_1183 & _GEN_1098 : ~_GEN_1130 & _GEN_1098;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1227 = _GEN_31 ? ~_GEN_1185 & _GEN_1099 : ~_GEN_1131 & _GEN_1099;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1228 = _GEN_31 ? ~_GEN_1187 & _GEN_1100 : ~_GEN_1132 & _GEN_1100;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1229 = _GEN_31 ? ~_GEN_1189 & _GEN_1101 : ~_GEN_1133 & _GEN_1101;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1230 = _GEN_31 ? ~_GEN_1191 & _GEN_1102 : ~_GEN_1134 & _GEN_1102;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1231 = _GEN_31 ? ~_GEN_1193 & _GEN_1103 : ~_GEN_1135 & _GEN_1103;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1232 = _GEN_31 ? ~_GEN_1195 & _GEN_1104 : ~_GEN_1136 & _GEN_1104;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1233 = _GEN_31 ? ~_GEN_1197 & _GEN_1105 : ~_GEN_1137 & _GEN_1105;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1234 = _GEN_31 ? ~_GEN_1199 & _GEN_1106 : ~_GEN_1138 & _GEN_1106;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1235 = _GEN_31 ? ~_GEN_1201 & _GEN_1107 : ~_GEN_1139 & _GEN_1107;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1236 = _GEN_31 ? ~_GEN_1203 & _GEN_1108 : ~_GEN_1140 & _GEN_1108;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1270 = _GEN_33 ? ~_GEN_1269 & _GEN_1142 : ~_GEN_1237 & _GEN_1142;	// rob.scala:346:{27,69}, :347:31
    _GEN_1272 = _GEN_33 ? ~_GEN_1271 & _GEN_1144 : ~_GEN_1238 & _GEN_1144;	// rob.scala:346:{27,69}, :347:31
    _GEN_1274 = _GEN_33 ? ~_GEN_1273 & _GEN_1146 : ~_GEN_1239 & _GEN_1146;	// rob.scala:346:{27,69}, :347:31
    _GEN_1276 = _GEN_33 ? ~_GEN_1275 & _GEN_1148 : ~_GEN_1240 & _GEN_1148;	// rob.scala:346:{27,69}, :347:31
    _GEN_1278 = _GEN_33 ? ~_GEN_1277 & _GEN_1150 : ~_GEN_1241 & _GEN_1150;	// rob.scala:346:{27,69}, :347:31
    _GEN_1280 = _GEN_33 ? ~_GEN_1279 & _GEN_1152 : ~_GEN_1242 & _GEN_1152;	// rob.scala:346:{27,69}, :347:31
    _GEN_1282 = _GEN_33 ? ~_GEN_1281 & _GEN_1154 : ~_GEN_1243 & _GEN_1154;	// rob.scala:346:{27,69}, :347:31
    _GEN_1284 = _GEN_33 ? ~_GEN_1283 & _GEN_1156 : ~_GEN_1244 & _GEN_1156;	// rob.scala:346:{27,69}, :347:31
    _GEN_1286 = _GEN_33 ? ~_GEN_1285 & _GEN_1158 : ~_GEN_1245 & _GEN_1158;	// rob.scala:346:{27,69}, :347:31
    _GEN_1288 = _GEN_33 ? ~_GEN_1287 & _GEN_1160 : ~_GEN_1246 & _GEN_1160;	// rob.scala:346:{27,69}, :347:31
    _GEN_1290 = _GEN_33 ? ~_GEN_1289 & _GEN_1162 : ~_GEN_1247 & _GEN_1162;	// rob.scala:346:{27,69}, :347:31
    _GEN_1292 = _GEN_33 ? ~_GEN_1291 & _GEN_1164 : ~_GEN_1248 & _GEN_1164;	// rob.scala:346:{27,69}, :347:31
    _GEN_1294 = _GEN_33 ? ~_GEN_1293 & _GEN_1166 : ~_GEN_1249 & _GEN_1166;	// rob.scala:346:{27,69}, :347:31
    _GEN_1296 = _GEN_33 ? ~_GEN_1295 & _GEN_1168 : ~_GEN_1250 & _GEN_1168;	// rob.scala:346:{27,69}, :347:31
    _GEN_1298 = _GEN_33 ? ~_GEN_1297 & _GEN_1170 : ~_GEN_1251 & _GEN_1170;	// rob.scala:346:{27,69}, :347:31
    _GEN_1300 = _GEN_33 ? ~_GEN_1299 & _GEN_1172 : ~_GEN_1252 & _GEN_1172;	// rob.scala:346:{27,69}, :347:31
    _GEN_1302 = _GEN_33 ? ~_GEN_1301 & _GEN_1174 : ~_GEN_1253 & _GEN_1174;	// rob.scala:346:{27,69}, :347:31
    _GEN_1304 = _GEN_33 ? ~_GEN_1303 & _GEN_1176 : ~_GEN_1254 & _GEN_1176;	// rob.scala:346:{27,69}, :347:31
    _GEN_1306 = _GEN_33 ? ~_GEN_1305 & _GEN_1178 : ~_GEN_1255 & _GEN_1178;	// rob.scala:346:{27,69}, :347:31
    _GEN_1308 = _GEN_33 ? ~_GEN_1307 & _GEN_1180 : ~_GEN_1256 & _GEN_1180;	// rob.scala:346:{27,69}, :347:31
    _GEN_1310 = _GEN_33 ? ~_GEN_1309 & _GEN_1182 : ~_GEN_1257 & _GEN_1182;	// rob.scala:346:{27,69}, :347:31
    _GEN_1312 = _GEN_33 ? ~_GEN_1311 & _GEN_1184 : ~_GEN_1258 & _GEN_1184;	// rob.scala:346:{27,69}, :347:31
    _GEN_1314 = _GEN_33 ? ~_GEN_1313 & _GEN_1186 : ~_GEN_1259 & _GEN_1186;	// rob.scala:346:{27,69}, :347:31
    _GEN_1316 = _GEN_33 ? ~_GEN_1315 & _GEN_1188 : ~_GEN_1260 & _GEN_1188;	// rob.scala:346:{27,69}, :347:31
    _GEN_1318 = _GEN_33 ? ~_GEN_1317 & _GEN_1190 : ~_GEN_1261 & _GEN_1190;	// rob.scala:346:{27,69}, :347:31
    _GEN_1320 = _GEN_33 ? ~_GEN_1319 & _GEN_1192 : ~_GEN_1262 & _GEN_1192;	// rob.scala:346:{27,69}, :347:31
    _GEN_1322 = _GEN_33 ? ~_GEN_1321 & _GEN_1194 : ~_GEN_1263 & _GEN_1194;	// rob.scala:346:{27,69}, :347:31
    _GEN_1324 = _GEN_33 ? ~_GEN_1323 & _GEN_1196 : ~_GEN_1264 & _GEN_1196;	// rob.scala:346:{27,69}, :347:31
    _GEN_1326 = _GEN_33 ? ~_GEN_1325 & _GEN_1198 : ~_GEN_1265 & _GEN_1198;	// rob.scala:346:{27,69}, :347:31
    _GEN_1328 = _GEN_33 ? ~_GEN_1327 & _GEN_1200 : ~_GEN_1266 & _GEN_1200;	// rob.scala:346:{27,69}, :347:31
    _GEN_1330 = _GEN_33 ? ~_GEN_1329 & _GEN_1202 : ~_GEN_1267 & _GEN_1202;	// rob.scala:346:{27,69}, :347:31
    _GEN_1332 = _GEN_33 ? ~_GEN_1331 & _GEN_1204 : ~_GEN_1268 & _GEN_1204;	// rob.scala:346:{27,69}, :347:31
    _GEN_1333 = _GEN_33 ? ~_GEN_1269 & _GEN_1205 : ~_GEN_1237 & _GEN_1205;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1334 = _GEN_33 ? ~_GEN_1271 & _GEN_1206 : ~_GEN_1238 & _GEN_1206;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1335 = _GEN_33 ? ~_GEN_1273 & _GEN_1207 : ~_GEN_1239 & _GEN_1207;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1336 = _GEN_33 ? ~_GEN_1275 & _GEN_1208 : ~_GEN_1240 & _GEN_1208;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1337 = _GEN_33 ? ~_GEN_1277 & _GEN_1209 : ~_GEN_1241 & _GEN_1209;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1338 = _GEN_33 ? ~_GEN_1279 & _GEN_1210 : ~_GEN_1242 & _GEN_1210;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1339 = _GEN_33 ? ~_GEN_1281 & _GEN_1211 : ~_GEN_1243 & _GEN_1211;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1340 = _GEN_33 ? ~_GEN_1283 & _GEN_1212 : ~_GEN_1244 & _GEN_1212;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1341 = _GEN_33 ? ~_GEN_1285 & _GEN_1213 : ~_GEN_1245 & _GEN_1213;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1342 = _GEN_33 ? ~_GEN_1287 & _GEN_1214 : ~_GEN_1246 & _GEN_1214;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1343 = _GEN_33 ? ~_GEN_1289 & _GEN_1215 : ~_GEN_1247 & _GEN_1215;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1344 = _GEN_33 ? ~_GEN_1291 & _GEN_1216 : ~_GEN_1248 & _GEN_1216;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1345 = _GEN_33 ? ~_GEN_1293 & _GEN_1217 : ~_GEN_1249 & _GEN_1217;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1346 = _GEN_33 ? ~_GEN_1295 & _GEN_1218 : ~_GEN_1250 & _GEN_1218;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1347 = _GEN_33 ? ~_GEN_1297 & _GEN_1219 : ~_GEN_1251 & _GEN_1219;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1348 = _GEN_33 ? ~_GEN_1299 & _GEN_1220 : ~_GEN_1252 & _GEN_1220;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1349 = _GEN_33 ? ~_GEN_1301 & _GEN_1221 : ~_GEN_1253 & _GEN_1221;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1350 = _GEN_33 ? ~_GEN_1303 & _GEN_1222 : ~_GEN_1254 & _GEN_1222;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1351 = _GEN_33 ? ~_GEN_1305 & _GEN_1223 : ~_GEN_1255 & _GEN_1223;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1352 = _GEN_33 ? ~_GEN_1307 & _GEN_1224 : ~_GEN_1256 & _GEN_1224;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1353 = _GEN_33 ? ~_GEN_1309 & _GEN_1225 : ~_GEN_1257 & _GEN_1225;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1354 = _GEN_33 ? ~_GEN_1311 & _GEN_1226 : ~_GEN_1258 & _GEN_1226;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1355 = _GEN_33 ? ~_GEN_1313 & _GEN_1227 : ~_GEN_1259 & _GEN_1227;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1356 = _GEN_33 ? ~_GEN_1315 & _GEN_1228 : ~_GEN_1260 & _GEN_1228;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1357 = _GEN_33 ? ~_GEN_1317 & _GEN_1229 : ~_GEN_1261 & _GEN_1229;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1358 = _GEN_33 ? ~_GEN_1319 & _GEN_1230 : ~_GEN_1262 & _GEN_1230;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1359 = _GEN_33 ? ~_GEN_1321 & _GEN_1231 : ~_GEN_1263 & _GEN_1231;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1360 = _GEN_33 ? ~_GEN_1323 & _GEN_1232 : ~_GEN_1264 & _GEN_1232;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1361 = _GEN_33 ? ~_GEN_1325 & _GEN_1233 : ~_GEN_1265 & _GEN_1233;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1362 = _GEN_33 ? ~_GEN_1327 & _GEN_1234 : ~_GEN_1266 & _GEN_1234;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1363 = _GEN_33 ? ~_GEN_1329 & _GEN_1235 : ~_GEN_1267 & _GEN_1235;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1364 = _GEN_33 ? ~_GEN_1331 & _GEN_1236 : ~_GEN_1268 & _GEN_1236;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1398 = _GEN_35 ? ~_GEN_1397 & _GEN_1270 : ~_GEN_1365 & _GEN_1270;	// rob.scala:346:{27,69}, :347:31
    _GEN_1400 = _GEN_35 ? ~_GEN_1399 & _GEN_1272 : ~_GEN_1366 & _GEN_1272;	// rob.scala:346:{27,69}, :347:31
    _GEN_1402 = _GEN_35 ? ~_GEN_1401 & _GEN_1274 : ~_GEN_1367 & _GEN_1274;	// rob.scala:346:{27,69}, :347:31
    _GEN_1404 = _GEN_35 ? ~_GEN_1403 & _GEN_1276 : ~_GEN_1368 & _GEN_1276;	// rob.scala:346:{27,69}, :347:31
    _GEN_1406 = _GEN_35 ? ~_GEN_1405 & _GEN_1278 : ~_GEN_1369 & _GEN_1278;	// rob.scala:346:{27,69}, :347:31
    _GEN_1408 = _GEN_35 ? ~_GEN_1407 & _GEN_1280 : ~_GEN_1370 & _GEN_1280;	// rob.scala:346:{27,69}, :347:31
    _GEN_1410 = _GEN_35 ? ~_GEN_1409 & _GEN_1282 : ~_GEN_1371 & _GEN_1282;	// rob.scala:346:{27,69}, :347:31
    _GEN_1412 = _GEN_35 ? ~_GEN_1411 & _GEN_1284 : ~_GEN_1372 & _GEN_1284;	// rob.scala:346:{27,69}, :347:31
    _GEN_1414 = _GEN_35 ? ~_GEN_1413 & _GEN_1286 : ~_GEN_1373 & _GEN_1286;	// rob.scala:346:{27,69}, :347:31
    _GEN_1416 = _GEN_35 ? ~_GEN_1415 & _GEN_1288 : ~_GEN_1374 & _GEN_1288;	// rob.scala:346:{27,69}, :347:31
    _GEN_1418 = _GEN_35 ? ~_GEN_1417 & _GEN_1290 : ~_GEN_1375 & _GEN_1290;	// rob.scala:346:{27,69}, :347:31
    _GEN_1420 = _GEN_35 ? ~_GEN_1419 & _GEN_1292 : ~_GEN_1376 & _GEN_1292;	// rob.scala:346:{27,69}, :347:31
    _GEN_1422 = _GEN_35 ? ~_GEN_1421 & _GEN_1294 : ~_GEN_1377 & _GEN_1294;	// rob.scala:346:{27,69}, :347:31
    _GEN_1424 = _GEN_35 ? ~_GEN_1423 & _GEN_1296 : ~_GEN_1378 & _GEN_1296;	// rob.scala:346:{27,69}, :347:31
    _GEN_1426 = _GEN_35 ? ~_GEN_1425 & _GEN_1298 : ~_GEN_1379 & _GEN_1298;	// rob.scala:346:{27,69}, :347:31
    _GEN_1428 = _GEN_35 ? ~_GEN_1427 & _GEN_1300 : ~_GEN_1380 & _GEN_1300;	// rob.scala:346:{27,69}, :347:31
    _GEN_1430 = _GEN_35 ? ~_GEN_1429 & _GEN_1302 : ~_GEN_1381 & _GEN_1302;	// rob.scala:346:{27,69}, :347:31
    _GEN_1432 = _GEN_35 ? ~_GEN_1431 & _GEN_1304 : ~_GEN_1382 & _GEN_1304;	// rob.scala:346:{27,69}, :347:31
    _GEN_1434 = _GEN_35 ? ~_GEN_1433 & _GEN_1306 : ~_GEN_1383 & _GEN_1306;	// rob.scala:346:{27,69}, :347:31
    _GEN_1436 = _GEN_35 ? ~_GEN_1435 & _GEN_1308 : ~_GEN_1384 & _GEN_1308;	// rob.scala:346:{27,69}, :347:31
    _GEN_1438 = _GEN_35 ? ~_GEN_1437 & _GEN_1310 : ~_GEN_1385 & _GEN_1310;	// rob.scala:346:{27,69}, :347:31
    _GEN_1440 = _GEN_35 ? ~_GEN_1439 & _GEN_1312 : ~_GEN_1386 & _GEN_1312;	// rob.scala:346:{27,69}, :347:31
    _GEN_1442 = _GEN_35 ? ~_GEN_1441 & _GEN_1314 : ~_GEN_1387 & _GEN_1314;	// rob.scala:346:{27,69}, :347:31
    _GEN_1444 = _GEN_35 ? ~_GEN_1443 & _GEN_1316 : ~_GEN_1388 & _GEN_1316;	// rob.scala:346:{27,69}, :347:31
    _GEN_1446 = _GEN_35 ? ~_GEN_1445 & _GEN_1318 : ~_GEN_1389 & _GEN_1318;	// rob.scala:346:{27,69}, :347:31
    _GEN_1448 = _GEN_35 ? ~_GEN_1447 & _GEN_1320 : ~_GEN_1390 & _GEN_1320;	// rob.scala:346:{27,69}, :347:31
    _GEN_1450 = _GEN_35 ? ~_GEN_1449 & _GEN_1322 : ~_GEN_1391 & _GEN_1322;	// rob.scala:346:{27,69}, :347:31
    _GEN_1452 = _GEN_35 ? ~_GEN_1451 & _GEN_1324 : ~_GEN_1392 & _GEN_1324;	// rob.scala:346:{27,69}, :347:31
    _GEN_1454 = _GEN_35 ? ~_GEN_1453 & _GEN_1326 : ~_GEN_1393 & _GEN_1326;	// rob.scala:346:{27,69}, :347:31
    _GEN_1456 = _GEN_35 ? ~_GEN_1455 & _GEN_1328 : ~_GEN_1394 & _GEN_1328;	// rob.scala:346:{27,69}, :347:31
    _GEN_1458 = _GEN_35 ? ~_GEN_1457 & _GEN_1330 : ~_GEN_1395 & _GEN_1330;	// rob.scala:346:{27,69}, :347:31
    _GEN_1460 = _GEN_35 ? ~_GEN_1459 & _GEN_1332 : ~_GEN_1396 & _GEN_1332;	// rob.scala:346:{27,69}, :347:31
    _GEN_1461 = _GEN_35 ? ~_GEN_1397 & _GEN_1333 : ~_GEN_1365 & _GEN_1333;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1462 = _GEN_35 ? ~_GEN_1399 & _GEN_1334 : ~_GEN_1366 & _GEN_1334;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1463 = _GEN_35 ? ~_GEN_1401 & _GEN_1335 : ~_GEN_1367 & _GEN_1335;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1464 = _GEN_35 ? ~_GEN_1403 & _GEN_1336 : ~_GEN_1368 & _GEN_1336;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1465 = _GEN_35 ? ~_GEN_1405 & _GEN_1337 : ~_GEN_1369 & _GEN_1337;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1466 = _GEN_35 ? ~_GEN_1407 & _GEN_1338 : ~_GEN_1370 & _GEN_1338;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1467 = _GEN_35 ? ~_GEN_1409 & _GEN_1339 : ~_GEN_1371 & _GEN_1339;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1468 = _GEN_35 ? ~_GEN_1411 & _GEN_1340 : ~_GEN_1372 & _GEN_1340;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1469 = _GEN_35 ? ~_GEN_1413 & _GEN_1341 : ~_GEN_1373 & _GEN_1341;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1470 = _GEN_35 ? ~_GEN_1415 & _GEN_1342 : ~_GEN_1374 & _GEN_1342;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1471 = _GEN_35 ? ~_GEN_1417 & _GEN_1343 : ~_GEN_1375 & _GEN_1343;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1472 = _GEN_35 ? ~_GEN_1419 & _GEN_1344 : ~_GEN_1376 & _GEN_1344;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1473 = _GEN_35 ? ~_GEN_1421 & _GEN_1345 : ~_GEN_1377 & _GEN_1345;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1474 = _GEN_35 ? ~_GEN_1423 & _GEN_1346 : ~_GEN_1378 & _GEN_1346;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1475 = _GEN_35 ? ~_GEN_1425 & _GEN_1347 : ~_GEN_1379 & _GEN_1347;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1476 = _GEN_35 ? ~_GEN_1427 & _GEN_1348 : ~_GEN_1380 & _GEN_1348;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1477 = _GEN_35 ? ~_GEN_1429 & _GEN_1349 : ~_GEN_1381 & _GEN_1349;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1478 = _GEN_35 ? ~_GEN_1431 & _GEN_1350 : ~_GEN_1382 & _GEN_1350;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1479 = _GEN_35 ? ~_GEN_1433 & _GEN_1351 : ~_GEN_1383 & _GEN_1351;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1480 = _GEN_35 ? ~_GEN_1435 & _GEN_1352 : ~_GEN_1384 & _GEN_1352;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1481 = _GEN_35 ? ~_GEN_1437 & _GEN_1353 : ~_GEN_1385 & _GEN_1353;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1482 = _GEN_35 ? ~_GEN_1439 & _GEN_1354 : ~_GEN_1386 & _GEN_1354;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1483 = _GEN_35 ? ~_GEN_1441 & _GEN_1355 : ~_GEN_1387 & _GEN_1355;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1484 = _GEN_35 ? ~_GEN_1443 & _GEN_1356 : ~_GEN_1388 & _GEN_1356;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1485 = _GEN_35 ? ~_GEN_1445 & _GEN_1357 : ~_GEN_1389 & _GEN_1357;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1486 = _GEN_35 ? ~_GEN_1447 & _GEN_1358 : ~_GEN_1390 & _GEN_1358;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1487 = _GEN_35 ? ~_GEN_1449 & _GEN_1359 : ~_GEN_1391 & _GEN_1359;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1488 = _GEN_35 ? ~_GEN_1451 & _GEN_1360 : ~_GEN_1392 & _GEN_1360;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1489 = _GEN_35 ? ~_GEN_1453 & _GEN_1361 : ~_GEN_1393 & _GEN_1361;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1490 = _GEN_35 ? ~_GEN_1455 & _GEN_1362 : ~_GEN_1394 & _GEN_1362;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1491 = _GEN_35 ? ~_GEN_1457 & _GEN_1363 : ~_GEN_1395 & _GEN_1363;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1492 = _GEN_35 ? ~_GEN_1459 & _GEN_1364 : ~_GEN_1396 & _GEN_1364;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1493 = _GEN_36 & _GEN_793;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1494 = _GEN_36 & _GEN_795;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1495 = _GEN_36 & _GEN_797;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1496 = _GEN_36 & _GEN_799;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1497 = _GEN_36 & _GEN_801;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1498 = _GEN_36 & _GEN_803;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1499 = _GEN_36 & _GEN_805;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1500 = _GEN_36 & _GEN_807;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1501 = _GEN_36 & _GEN_809;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1502 = _GEN_36 & _GEN_811;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1503 = _GEN_36 & _GEN_813;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1504 = _GEN_36 & _GEN_815;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1505 = _GEN_36 & _GEN_817;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1506 = _GEN_36 & _GEN_819;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1507 = _GEN_36 & _GEN_821;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1508 = _GEN_36 & _GEN_823;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1509 = _GEN_36 & _GEN_825;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1510 = _GEN_36 & _GEN_827;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1511 = _GEN_36 & _GEN_829;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1512 = _GEN_36 & _GEN_831;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1513 = _GEN_36 & _GEN_833;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1514 = _GEN_36 & _GEN_835;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1515 = _GEN_36 & _GEN_837;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1516 = _GEN_36 & _GEN_839;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1517 = _GEN_36 & _GEN_841;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1518 = _GEN_36 & _GEN_843;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1519 = _GEN_36 & _GEN_845;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1520 = _GEN_36 & _GEN_847;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1521 = _GEN_36 & _GEN_849;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1522 = _GEN_36 & _GEN_851;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1523 = _GEN_36 & _GEN_853;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_1524 = _GEN_36 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    _GEN_1525 = rbk_row_1 & _GEN_918;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1526 = rbk_row_1 & _GEN_920;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1527 = rbk_row_1 & _GEN_922;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1528 = rbk_row_1 & _GEN_924;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1529 = rbk_row_1 & _GEN_926;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1530 = rbk_row_1 & _GEN_928;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1531 = rbk_row_1 & _GEN_930;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1532 = rbk_row_1 & _GEN_932;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1533 = rbk_row_1 & _GEN_934;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1534 = rbk_row_1 & _GEN_936;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1535 = rbk_row_1 & _GEN_938;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1536 = rbk_row_1 & _GEN_940;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1537 = rbk_row_1 & _GEN_942;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1538 = rbk_row_1 & _GEN_944;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1539 = rbk_row_1 & _GEN_946;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1540 = rbk_row_1 & _GEN_948;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1541 = rbk_row_1 & _GEN_950;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1542 = rbk_row_1 & _GEN_952;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1543 = rbk_row_1 & _GEN_954;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1544 = rbk_row_1 & _GEN_956;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1545 = rbk_row_1 & _GEN_958;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1546 = rbk_row_1 & _GEN_960;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1547 = rbk_row_1 & _GEN_962;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1548 = rbk_row_1 & _GEN_964;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1549 = rbk_row_1 & _GEN_966;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1550 = rbk_row_1 & _GEN_968;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1551 = rbk_row_1 & _GEN_970;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1552 = rbk_row_1 & _GEN_972;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1553 = rbk_row_1 & _GEN_974;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1554 = rbk_row_1 & _GEN_976;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1555 = rbk_row_1 & _GEN_978;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_1556 = rbk_row_1 & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_1557 = io_brupdate_b1_mispredict_mask & rob_uop_1_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1558 = io_brupdate_b1_mispredict_mask & rob_uop_1_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1559 = io_brupdate_b1_mispredict_mask & rob_uop_1_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1560 = io_brupdate_b1_mispredict_mask & rob_uop_1_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1561 = io_brupdate_b1_mispredict_mask & rob_uop_1_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1562 = io_brupdate_b1_mispredict_mask & rob_uop_1_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1563 = io_brupdate_b1_mispredict_mask & rob_uop_1_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1564 = io_brupdate_b1_mispredict_mask & rob_uop_1_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1565 = io_brupdate_b1_mispredict_mask & rob_uop_1_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1566 = io_brupdate_b1_mispredict_mask & rob_uop_1_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1567 = io_brupdate_b1_mispredict_mask & rob_uop_1_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1568 = io_brupdate_b1_mispredict_mask & rob_uop_1_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1569 = io_brupdate_b1_mispredict_mask & rob_uop_1_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1570 = io_brupdate_b1_mispredict_mask & rob_uop_1_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1571 = io_brupdate_b1_mispredict_mask & rob_uop_1_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1572 = io_brupdate_b1_mispredict_mask & rob_uop_1_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1573 = io_brupdate_b1_mispredict_mask & rob_uop_1_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1574 = io_brupdate_b1_mispredict_mask & rob_uop_1_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1575 = io_brupdate_b1_mispredict_mask & rob_uop_1_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1576 = io_brupdate_b1_mispredict_mask & rob_uop_1_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1577 = io_brupdate_b1_mispredict_mask & rob_uop_1_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1578 = io_brupdate_b1_mispredict_mask & rob_uop_1_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1579 = io_brupdate_b1_mispredict_mask & rob_uop_1_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1580 = io_brupdate_b1_mispredict_mask & rob_uop_1_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1581 = io_brupdate_b1_mispredict_mask & rob_uop_1_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1582 = io_brupdate_b1_mispredict_mask & rob_uop_1_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1583 = io_brupdate_b1_mispredict_mask & rob_uop_1_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1584 = io_brupdate_b1_mispredict_mask & rob_uop_1_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1585 = io_brupdate_b1_mispredict_mask & rob_uop_1_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1586 = io_brupdate_b1_mispredict_mask & rob_uop_1_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1587 = io_brupdate_b1_mispredict_mask & rob_uop_1_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1588 = io_brupdate_b1_mispredict_mask & rob_uop_1_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_1589 = io_enq_valids_2 & _GEN_96;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1590 = io_enq_valids_2 & _GEN_98;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1591 = io_enq_valids_2 & _GEN_100;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1592 = io_enq_valids_2 & _GEN_102;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1593 = io_enq_valids_2 & _GEN_104;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1594 = io_enq_valids_2 & _GEN_106;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1595 = io_enq_valids_2 & _GEN_108;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1596 = io_enq_valids_2 & _GEN_110;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1597 = io_enq_valids_2 & _GEN_112;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1598 = io_enq_valids_2 & _GEN_114;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1599 = io_enq_valids_2 & _GEN_116;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1600 = io_enq_valids_2 & _GEN_118;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1601 = io_enq_valids_2 & _GEN_120;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1602 = io_enq_valids_2 & _GEN_122;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1603 = io_enq_valids_2 & _GEN_124;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1604 = io_enq_valids_2 & _GEN_126;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1605 = io_enq_valids_2 & _GEN_128;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1606 = io_enq_valids_2 & _GEN_130;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1607 = io_enq_valids_2 & _GEN_132;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1608 = io_enq_valids_2 & _GEN_134;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1609 = io_enq_valids_2 & _GEN_136;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1610 = io_enq_valids_2 & _GEN_138;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1611 = io_enq_valids_2 & _GEN_140;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1612 = io_enq_valids_2 & _GEN_142;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1613 = io_enq_valids_2 & _GEN_144;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1614 = io_enq_valids_2 & _GEN_146;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1615 = io_enq_valids_2 & _GEN_148;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1616 = io_enq_valids_2 & _GEN_150;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1617 = io_enq_valids_2 & _GEN_152;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1618 = io_enq_valids_2 & _GEN_154;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1619 = io_enq_valids_2 & _GEN_156;	// rob.scala:307:32, :323:29, :324:31
    _GEN_1620 = io_enq_valids_2 & (&rob_tail);	// rob.scala:228:29, :307:32, :323:29, :324:31
    _GEN_1621 = _GEN_1589 ? ~_rob_bsy_T_4 : rob_bsy_2_0;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1622 = _GEN_1590 ? ~_rob_bsy_T_4 : rob_bsy_2_1;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1623 = _GEN_1591 ? ~_rob_bsy_T_4 : rob_bsy_2_2;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1624 = _GEN_1592 ? ~_rob_bsy_T_4 : rob_bsy_2_3;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1625 = _GEN_1593 ? ~_rob_bsy_T_4 : rob_bsy_2_4;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1626 = _GEN_1594 ? ~_rob_bsy_T_4 : rob_bsy_2_5;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1627 = _GEN_1595 ? ~_rob_bsy_T_4 : rob_bsy_2_6;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1628 = _GEN_1596 ? ~_rob_bsy_T_4 : rob_bsy_2_7;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1629 = _GEN_1597 ? ~_rob_bsy_T_4 : rob_bsy_2_8;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1630 = _GEN_1598 ? ~_rob_bsy_T_4 : rob_bsy_2_9;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1631 = _GEN_1599 ? ~_rob_bsy_T_4 : rob_bsy_2_10;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1632 = _GEN_1600 ? ~_rob_bsy_T_4 : rob_bsy_2_11;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1633 = _GEN_1601 ? ~_rob_bsy_T_4 : rob_bsy_2_12;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1634 = _GEN_1602 ? ~_rob_bsy_T_4 : rob_bsy_2_13;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1635 = _GEN_1603 ? ~_rob_bsy_T_4 : rob_bsy_2_14;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1636 = _GEN_1604 ? ~_rob_bsy_T_4 : rob_bsy_2_15;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1637 = _GEN_1605 ? ~_rob_bsy_T_4 : rob_bsy_2_16;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1638 = _GEN_1606 ? ~_rob_bsy_T_4 : rob_bsy_2_17;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1639 = _GEN_1607 ? ~_rob_bsy_T_4 : rob_bsy_2_18;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1640 = _GEN_1608 ? ~_rob_bsy_T_4 : rob_bsy_2_19;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1641 = _GEN_1609 ? ~_rob_bsy_T_4 : rob_bsy_2_20;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1642 = _GEN_1610 ? ~_rob_bsy_T_4 : rob_bsy_2_21;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1643 = _GEN_1611 ? ~_rob_bsy_T_4 : rob_bsy_2_22;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1644 = _GEN_1612 ? ~_rob_bsy_T_4 : rob_bsy_2_23;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1645 = _GEN_1613 ? ~_rob_bsy_T_4 : rob_bsy_2_24;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1646 = _GEN_1614 ? ~_rob_bsy_T_4 : rob_bsy_2_25;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1647 = _GEN_1615 ? ~_rob_bsy_T_4 : rob_bsy_2_26;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1648 = _GEN_1616 ? ~_rob_bsy_T_4 : rob_bsy_2_27;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1649 = _GEN_1617 ? ~_rob_bsy_T_4 : rob_bsy_2_28;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1650 = _GEN_1618 ? ~_rob_bsy_T_4 : rob_bsy_2_29;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1651 = _GEN_1619 ? ~_rob_bsy_T_4 : rob_bsy_2_30;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1652 = _GEN_1620 ? ~_rob_bsy_T_4 : rob_bsy_2_31;	// rob.scala:307:32, :308:28, :323:29, :324:31, :325:{31,34,60}
    _GEN_1653 = _GEN_1589 ? _rob_unsafe_T_14 : rob_unsafe_2_0;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1654 = _GEN_1590 ? _rob_unsafe_T_14 : rob_unsafe_2_1;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1655 = _GEN_1591 ? _rob_unsafe_T_14 : rob_unsafe_2_2;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1656 = _GEN_1592 ? _rob_unsafe_T_14 : rob_unsafe_2_3;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1657 = _GEN_1593 ? _rob_unsafe_T_14 : rob_unsafe_2_4;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1658 = _GEN_1594 ? _rob_unsafe_T_14 : rob_unsafe_2_5;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1659 = _GEN_1595 ? _rob_unsafe_T_14 : rob_unsafe_2_6;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1660 = _GEN_1596 ? _rob_unsafe_T_14 : rob_unsafe_2_7;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1661 = _GEN_1597 ? _rob_unsafe_T_14 : rob_unsafe_2_8;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1662 = _GEN_1598 ? _rob_unsafe_T_14 : rob_unsafe_2_9;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1663 = _GEN_1599 ? _rob_unsafe_T_14 : rob_unsafe_2_10;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1664 = _GEN_1600 ? _rob_unsafe_T_14 : rob_unsafe_2_11;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1665 = _GEN_1601 ? _rob_unsafe_T_14 : rob_unsafe_2_12;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1666 = _GEN_1602 ? _rob_unsafe_T_14 : rob_unsafe_2_13;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1667 = _GEN_1603 ? _rob_unsafe_T_14 : rob_unsafe_2_14;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1668 = _GEN_1604 ? _rob_unsafe_T_14 : rob_unsafe_2_15;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1669 = _GEN_1605 ? _rob_unsafe_T_14 : rob_unsafe_2_16;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1670 = _GEN_1606 ? _rob_unsafe_T_14 : rob_unsafe_2_17;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1671 = _GEN_1607 ? _rob_unsafe_T_14 : rob_unsafe_2_18;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1672 = _GEN_1608 ? _rob_unsafe_T_14 : rob_unsafe_2_19;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1673 = _GEN_1609 ? _rob_unsafe_T_14 : rob_unsafe_2_20;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1674 = _GEN_1610 ? _rob_unsafe_T_14 : rob_unsafe_2_21;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1675 = _GEN_1611 ? _rob_unsafe_T_14 : rob_unsafe_2_22;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1676 = _GEN_1612 ? _rob_unsafe_T_14 : rob_unsafe_2_23;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1677 = _GEN_1613 ? _rob_unsafe_T_14 : rob_unsafe_2_24;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1678 = _GEN_1614 ? _rob_unsafe_T_14 : rob_unsafe_2_25;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1679 = _GEN_1615 ? _rob_unsafe_T_14 : rob_unsafe_2_26;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1680 = _GEN_1616 ? _rob_unsafe_T_14 : rob_unsafe_2_27;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1681 = _GEN_1617 ? _rob_unsafe_T_14 : rob_unsafe_2_28;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1682 = _GEN_1618 ? _rob_unsafe_T_14 : rob_unsafe_2_29;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1683 = _GEN_1619 ? _rob_unsafe_T_14 : rob_unsafe_2_30;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1684 = _GEN_1620 ? _rob_unsafe_T_14 : rob_unsafe_2_31;	// micro-op.scala:152:71, rob.scala:307:32, :309:28, :323:29, :324:31, :327:31
    _GEN_1718 = _GEN_61 ? ~_GEN_1717 & _GEN_1621 : ~_GEN_1685 & _GEN_1621;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1720 = _GEN_61 ? ~_GEN_1719 & _GEN_1622 : ~_GEN_1686 & _GEN_1622;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1722 = _GEN_61 ? ~_GEN_1721 & _GEN_1623 : ~_GEN_1687 & _GEN_1623;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1724 = _GEN_61 ? ~_GEN_1723 & _GEN_1624 : ~_GEN_1688 & _GEN_1624;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1726 = _GEN_61 ? ~_GEN_1725 & _GEN_1625 : ~_GEN_1689 & _GEN_1625;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1728 = _GEN_61 ? ~_GEN_1727 & _GEN_1626 : ~_GEN_1690 & _GEN_1626;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1730 = _GEN_61 ? ~_GEN_1729 & _GEN_1627 : ~_GEN_1691 & _GEN_1627;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1732 = _GEN_61 ? ~_GEN_1731 & _GEN_1628 : ~_GEN_1692 & _GEN_1628;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1734 = _GEN_61 ? ~_GEN_1733 & _GEN_1629 : ~_GEN_1693 & _GEN_1629;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1736 = _GEN_61 ? ~_GEN_1735 & _GEN_1630 : ~_GEN_1694 & _GEN_1630;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1738 = _GEN_61 ? ~_GEN_1737 & _GEN_1631 : ~_GEN_1695 & _GEN_1631;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1740 = _GEN_61 ? ~_GEN_1739 & _GEN_1632 : ~_GEN_1696 & _GEN_1632;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1742 = _GEN_61 ? ~_GEN_1741 & _GEN_1633 : ~_GEN_1697 & _GEN_1633;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1744 = _GEN_61 ? ~_GEN_1743 & _GEN_1634 : ~_GEN_1698 & _GEN_1634;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1746 = _GEN_61 ? ~_GEN_1745 & _GEN_1635 : ~_GEN_1699 & _GEN_1635;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1748 = _GEN_61 ? ~_GEN_1747 & _GEN_1636 : ~_GEN_1700 & _GEN_1636;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1750 = _GEN_61 ? ~_GEN_1749 & _GEN_1637 : ~_GEN_1701 & _GEN_1637;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1752 = _GEN_61 ? ~_GEN_1751 & _GEN_1638 : ~_GEN_1702 & _GEN_1638;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1754 = _GEN_61 ? ~_GEN_1753 & _GEN_1639 : ~_GEN_1703 & _GEN_1639;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1756 = _GEN_61 ? ~_GEN_1755 & _GEN_1640 : ~_GEN_1704 & _GEN_1640;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1758 = _GEN_61 ? ~_GEN_1757 & _GEN_1641 : ~_GEN_1705 & _GEN_1641;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1760 = _GEN_61 ? ~_GEN_1759 & _GEN_1642 : ~_GEN_1706 & _GEN_1642;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1762 = _GEN_61 ? ~_GEN_1761 & _GEN_1643 : ~_GEN_1707 & _GEN_1643;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1764 = _GEN_61 ? ~_GEN_1763 & _GEN_1644 : ~_GEN_1708 & _GEN_1644;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1766 = _GEN_61 ? ~_GEN_1765 & _GEN_1645 : ~_GEN_1709 & _GEN_1645;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1768 = _GEN_61 ? ~_GEN_1767 & _GEN_1646 : ~_GEN_1710 & _GEN_1646;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1770 = _GEN_61 ? ~_GEN_1769 & _GEN_1647 : ~_GEN_1711 & _GEN_1647;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1772 = _GEN_61 ? ~_GEN_1771 & _GEN_1648 : ~_GEN_1712 & _GEN_1648;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1774 = _GEN_61 ? ~_GEN_1773 & _GEN_1649 : ~_GEN_1713 & _GEN_1649;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1776 = _GEN_61 ? ~_GEN_1775 & _GEN_1650 : ~_GEN_1714 & _GEN_1650;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1778 = _GEN_61 ? ~_GEN_1777 & _GEN_1651 : ~_GEN_1715 & _GEN_1651;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1780 = _GEN_61 ? ~_GEN_1779 & _GEN_1652 : ~_GEN_1716 & _GEN_1652;	// rob.scala:308:28, :323:29, :325:31, :346:{27,69}, :347:31
    _GEN_1781 = _GEN_61 ? ~_GEN_1717 & _GEN_1653 : ~_GEN_1685 & _GEN_1653;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1782 = _GEN_61 ? ~_GEN_1719 & _GEN_1654 : ~_GEN_1686 & _GEN_1654;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1783 = _GEN_61 ? ~_GEN_1721 & _GEN_1655 : ~_GEN_1687 & _GEN_1655;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1784 = _GEN_61 ? ~_GEN_1723 & _GEN_1656 : ~_GEN_1688 & _GEN_1656;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1785 = _GEN_61 ? ~_GEN_1725 & _GEN_1657 : ~_GEN_1689 & _GEN_1657;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1786 = _GEN_61 ? ~_GEN_1727 & _GEN_1658 : ~_GEN_1690 & _GEN_1658;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1787 = _GEN_61 ? ~_GEN_1729 & _GEN_1659 : ~_GEN_1691 & _GEN_1659;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1788 = _GEN_61 ? ~_GEN_1731 & _GEN_1660 : ~_GEN_1692 & _GEN_1660;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1789 = _GEN_61 ? ~_GEN_1733 & _GEN_1661 : ~_GEN_1693 & _GEN_1661;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1790 = _GEN_61 ? ~_GEN_1735 & _GEN_1662 : ~_GEN_1694 & _GEN_1662;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1791 = _GEN_61 ? ~_GEN_1737 & _GEN_1663 : ~_GEN_1695 & _GEN_1663;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1792 = _GEN_61 ? ~_GEN_1739 & _GEN_1664 : ~_GEN_1696 & _GEN_1664;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1793 = _GEN_61 ? ~_GEN_1741 & _GEN_1665 : ~_GEN_1697 & _GEN_1665;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1794 = _GEN_61 ? ~_GEN_1743 & _GEN_1666 : ~_GEN_1698 & _GEN_1666;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1795 = _GEN_61 ? ~_GEN_1745 & _GEN_1667 : ~_GEN_1699 & _GEN_1667;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1796 = _GEN_61 ? ~_GEN_1747 & _GEN_1668 : ~_GEN_1700 & _GEN_1668;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1797 = _GEN_61 ? ~_GEN_1749 & _GEN_1669 : ~_GEN_1701 & _GEN_1669;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1798 = _GEN_61 ? ~_GEN_1751 & _GEN_1670 : ~_GEN_1702 & _GEN_1670;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1799 = _GEN_61 ? ~_GEN_1753 & _GEN_1671 : ~_GEN_1703 & _GEN_1671;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1800 = _GEN_61 ? ~_GEN_1755 & _GEN_1672 : ~_GEN_1704 & _GEN_1672;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1801 = _GEN_61 ? ~_GEN_1757 & _GEN_1673 : ~_GEN_1705 & _GEN_1673;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1802 = _GEN_61 ? ~_GEN_1759 & _GEN_1674 : ~_GEN_1706 & _GEN_1674;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1803 = _GEN_61 ? ~_GEN_1761 & _GEN_1675 : ~_GEN_1707 & _GEN_1675;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1804 = _GEN_61 ? ~_GEN_1763 & _GEN_1676 : ~_GEN_1708 & _GEN_1676;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1805 = _GEN_61 ? ~_GEN_1765 & _GEN_1677 : ~_GEN_1709 & _GEN_1677;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1806 = _GEN_61 ? ~_GEN_1767 & _GEN_1678 : ~_GEN_1710 & _GEN_1678;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1807 = _GEN_61 ? ~_GEN_1769 & _GEN_1679 : ~_GEN_1711 & _GEN_1679;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1808 = _GEN_61 ? ~_GEN_1771 & _GEN_1680 : ~_GEN_1712 & _GEN_1680;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1809 = _GEN_61 ? ~_GEN_1773 & _GEN_1681 : ~_GEN_1713 & _GEN_1681;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1810 = _GEN_61 ? ~_GEN_1775 & _GEN_1682 : ~_GEN_1714 & _GEN_1682;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1811 = _GEN_61 ? ~_GEN_1777 & _GEN_1683 : ~_GEN_1715 & _GEN_1683;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1812 = _GEN_61 ? ~_GEN_1779 & _GEN_1684 : ~_GEN_1716 & _GEN_1684;	// rob.scala:309:28, :323:29, :327:31, :346:{27,69}, :347:31, :348:31
    _GEN_1846 = _GEN_63 ? ~_GEN_1845 & _GEN_1718 : ~_GEN_1813 & _GEN_1718;	// rob.scala:346:{27,69}, :347:31
    _GEN_1848 = _GEN_63 ? ~_GEN_1847 & _GEN_1720 : ~_GEN_1814 & _GEN_1720;	// rob.scala:346:{27,69}, :347:31
    _GEN_1850 = _GEN_63 ? ~_GEN_1849 & _GEN_1722 : ~_GEN_1815 & _GEN_1722;	// rob.scala:346:{27,69}, :347:31
    _GEN_1852 = _GEN_63 ? ~_GEN_1851 & _GEN_1724 : ~_GEN_1816 & _GEN_1724;	// rob.scala:346:{27,69}, :347:31
    _GEN_1854 = _GEN_63 ? ~_GEN_1853 & _GEN_1726 : ~_GEN_1817 & _GEN_1726;	// rob.scala:346:{27,69}, :347:31
    _GEN_1856 = _GEN_63 ? ~_GEN_1855 & _GEN_1728 : ~_GEN_1818 & _GEN_1728;	// rob.scala:346:{27,69}, :347:31
    _GEN_1858 = _GEN_63 ? ~_GEN_1857 & _GEN_1730 : ~_GEN_1819 & _GEN_1730;	// rob.scala:346:{27,69}, :347:31
    _GEN_1860 = _GEN_63 ? ~_GEN_1859 & _GEN_1732 : ~_GEN_1820 & _GEN_1732;	// rob.scala:346:{27,69}, :347:31
    _GEN_1862 = _GEN_63 ? ~_GEN_1861 & _GEN_1734 : ~_GEN_1821 & _GEN_1734;	// rob.scala:346:{27,69}, :347:31
    _GEN_1864 = _GEN_63 ? ~_GEN_1863 & _GEN_1736 : ~_GEN_1822 & _GEN_1736;	// rob.scala:346:{27,69}, :347:31
    _GEN_1866 = _GEN_63 ? ~_GEN_1865 & _GEN_1738 : ~_GEN_1823 & _GEN_1738;	// rob.scala:346:{27,69}, :347:31
    _GEN_1868 = _GEN_63 ? ~_GEN_1867 & _GEN_1740 : ~_GEN_1824 & _GEN_1740;	// rob.scala:346:{27,69}, :347:31
    _GEN_1870 = _GEN_63 ? ~_GEN_1869 & _GEN_1742 : ~_GEN_1825 & _GEN_1742;	// rob.scala:346:{27,69}, :347:31
    _GEN_1872 = _GEN_63 ? ~_GEN_1871 & _GEN_1744 : ~_GEN_1826 & _GEN_1744;	// rob.scala:346:{27,69}, :347:31
    _GEN_1874 = _GEN_63 ? ~_GEN_1873 & _GEN_1746 : ~_GEN_1827 & _GEN_1746;	// rob.scala:346:{27,69}, :347:31
    _GEN_1876 = _GEN_63 ? ~_GEN_1875 & _GEN_1748 : ~_GEN_1828 & _GEN_1748;	// rob.scala:346:{27,69}, :347:31
    _GEN_1878 = _GEN_63 ? ~_GEN_1877 & _GEN_1750 : ~_GEN_1829 & _GEN_1750;	// rob.scala:346:{27,69}, :347:31
    _GEN_1880 = _GEN_63 ? ~_GEN_1879 & _GEN_1752 : ~_GEN_1830 & _GEN_1752;	// rob.scala:346:{27,69}, :347:31
    _GEN_1882 = _GEN_63 ? ~_GEN_1881 & _GEN_1754 : ~_GEN_1831 & _GEN_1754;	// rob.scala:346:{27,69}, :347:31
    _GEN_1884 = _GEN_63 ? ~_GEN_1883 & _GEN_1756 : ~_GEN_1832 & _GEN_1756;	// rob.scala:346:{27,69}, :347:31
    _GEN_1886 = _GEN_63 ? ~_GEN_1885 & _GEN_1758 : ~_GEN_1833 & _GEN_1758;	// rob.scala:346:{27,69}, :347:31
    _GEN_1888 = _GEN_63 ? ~_GEN_1887 & _GEN_1760 : ~_GEN_1834 & _GEN_1760;	// rob.scala:346:{27,69}, :347:31
    _GEN_1890 = _GEN_63 ? ~_GEN_1889 & _GEN_1762 : ~_GEN_1835 & _GEN_1762;	// rob.scala:346:{27,69}, :347:31
    _GEN_1892 = _GEN_63 ? ~_GEN_1891 & _GEN_1764 : ~_GEN_1836 & _GEN_1764;	// rob.scala:346:{27,69}, :347:31
    _GEN_1894 = _GEN_63 ? ~_GEN_1893 & _GEN_1766 : ~_GEN_1837 & _GEN_1766;	// rob.scala:346:{27,69}, :347:31
    _GEN_1896 = _GEN_63 ? ~_GEN_1895 & _GEN_1768 : ~_GEN_1838 & _GEN_1768;	// rob.scala:346:{27,69}, :347:31
    _GEN_1898 = _GEN_63 ? ~_GEN_1897 & _GEN_1770 : ~_GEN_1839 & _GEN_1770;	// rob.scala:346:{27,69}, :347:31
    _GEN_1900 = _GEN_63 ? ~_GEN_1899 & _GEN_1772 : ~_GEN_1840 & _GEN_1772;	// rob.scala:346:{27,69}, :347:31
    _GEN_1902 = _GEN_63 ? ~_GEN_1901 & _GEN_1774 : ~_GEN_1841 & _GEN_1774;	// rob.scala:346:{27,69}, :347:31
    _GEN_1904 = _GEN_63 ? ~_GEN_1903 & _GEN_1776 : ~_GEN_1842 & _GEN_1776;	// rob.scala:346:{27,69}, :347:31
    _GEN_1906 = _GEN_63 ? ~_GEN_1905 & _GEN_1778 : ~_GEN_1843 & _GEN_1778;	// rob.scala:346:{27,69}, :347:31
    _GEN_1908 = _GEN_63 ? ~_GEN_1907 & _GEN_1780 : ~_GEN_1844 & _GEN_1780;	// rob.scala:346:{27,69}, :347:31
    _GEN_1909 = _GEN_63 ? ~_GEN_1845 & _GEN_1781 : ~_GEN_1813 & _GEN_1781;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1910 = _GEN_63 ? ~_GEN_1847 & _GEN_1782 : ~_GEN_1814 & _GEN_1782;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1911 = _GEN_63 ? ~_GEN_1849 & _GEN_1783 : ~_GEN_1815 & _GEN_1783;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1912 = _GEN_63 ? ~_GEN_1851 & _GEN_1784 : ~_GEN_1816 & _GEN_1784;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1913 = _GEN_63 ? ~_GEN_1853 & _GEN_1785 : ~_GEN_1817 & _GEN_1785;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1914 = _GEN_63 ? ~_GEN_1855 & _GEN_1786 : ~_GEN_1818 & _GEN_1786;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1915 = _GEN_63 ? ~_GEN_1857 & _GEN_1787 : ~_GEN_1819 & _GEN_1787;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1916 = _GEN_63 ? ~_GEN_1859 & _GEN_1788 : ~_GEN_1820 & _GEN_1788;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1917 = _GEN_63 ? ~_GEN_1861 & _GEN_1789 : ~_GEN_1821 & _GEN_1789;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1918 = _GEN_63 ? ~_GEN_1863 & _GEN_1790 : ~_GEN_1822 & _GEN_1790;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1919 = _GEN_63 ? ~_GEN_1865 & _GEN_1791 : ~_GEN_1823 & _GEN_1791;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1920 = _GEN_63 ? ~_GEN_1867 & _GEN_1792 : ~_GEN_1824 & _GEN_1792;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1921 = _GEN_63 ? ~_GEN_1869 & _GEN_1793 : ~_GEN_1825 & _GEN_1793;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1922 = _GEN_63 ? ~_GEN_1871 & _GEN_1794 : ~_GEN_1826 & _GEN_1794;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1923 = _GEN_63 ? ~_GEN_1873 & _GEN_1795 : ~_GEN_1827 & _GEN_1795;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1924 = _GEN_63 ? ~_GEN_1875 & _GEN_1796 : ~_GEN_1828 & _GEN_1796;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1925 = _GEN_63 ? ~_GEN_1877 & _GEN_1797 : ~_GEN_1829 & _GEN_1797;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1926 = _GEN_63 ? ~_GEN_1879 & _GEN_1798 : ~_GEN_1830 & _GEN_1798;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1927 = _GEN_63 ? ~_GEN_1881 & _GEN_1799 : ~_GEN_1831 & _GEN_1799;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1928 = _GEN_63 ? ~_GEN_1883 & _GEN_1800 : ~_GEN_1832 & _GEN_1800;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1929 = _GEN_63 ? ~_GEN_1885 & _GEN_1801 : ~_GEN_1833 & _GEN_1801;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1930 = _GEN_63 ? ~_GEN_1887 & _GEN_1802 : ~_GEN_1834 & _GEN_1802;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1931 = _GEN_63 ? ~_GEN_1889 & _GEN_1803 : ~_GEN_1835 & _GEN_1803;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1932 = _GEN_63 ? ~_GEN_1891 & _GEN_1804 : ~_GEN_1836 & _GEN_1804;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1933 = _GEN_63 ? ~_GEN_1893 & _GEN_1805 : ~_GEN_1837 & _GEN_1805;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1934 = _GEN_63 ? ~_GEN_1895 & _GEN_1806 : ~_GEN_1838 & _GEN_1806;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1935 = _GEN_63 ? ~_GEN_1897 & _GEN_1807 : ~_GEN_1839 & _GEN_1807;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1936 = _GEN_63 ? ~_GEN_1899 & _GEN_1808 : ~_GEN_1840 & _GEN_1808;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1937 = _GEN_63 ? ~_GEN_1901 & _GEN_1809 : ~_GEN_1841 & _GEN_1809;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1938 = _GEN_63 ? ~_GEN_1903 & _GEN_1810 : ~_GEN_1842 & _GEN_1810;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1939 = _GEN_63 ? ~_GEN_1905 & _GEN_1811 : ~_GEN_1843 & _GEN_1811;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1940 = _GEN_63 ? ~_GEN_1907 & _GEN_1812 : ~_GEN_1844 & _GEN_1812;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_1974 = _GEN_65 ? ~_GEN_1973 & _GEN_1846 : ~_GEN_1941 & _GEN_1846;	// rob.scala:346:{27,69}, :347:31
    _GEN_1976 = _GEN_65 ? ~_GEN_1975 & _GEN_1848 : ~_GEN_1942 & _GEN_1848;	// rob.scala:346:{27,69}, :347:31
    _GEN_1978 = _GEN_65 ? ~_GEN_1977 & _GEN_1850 : ~_GEN_1943 & _GEN_1850;	// rob.scala:346:{27,69}, :347:31
    _GEN_1980 = _GEN_65 ? ~_GEN_1979 & _GEN_1852 : ~_GEN_1944 & _GEN_1852;	// rob.scala:346:{27,69}, :347:31
    _GEN_1982 = _GEN_65 ? ~_GEN_1981 & _GEN_1854 : ~_GEN_1945 & _GEN_1854;	// rob.scala:346:{27,69}, :347:31
    _GEN_1984 = _GEN_65 ? ~_GEN_1983 & _GEN_1856 : ~_GEN_1946 & _GEN_1856;	// rob.scala:346:{27,69}, :347:31
    _GEN_1986 = _GEN_65 ? ~_GEN_1985 & _GEN_1858 : ~_GEN_1947 & _GEN_1858;	// rob.scala:346:{27,69}, :347:31
    _GEN_1988 = _GEN_65 ? ~_GEN_1987 & _GEN_1860 : ~_GEN_1948 & _GEN_1860;	// rob.scala:346:{27,69}, :347:31
    _GEN_1990 = _GEN_65 ? ~_GEN_1989 & _GEN_1862 : ~_GEN_1949 & _GEN_1862;	// rob.scala:346:{27,69}, :347:31
    _GEN_1992 = _GEN_65 ? ~_GEN_1991 & _GEN_1864 : ~_GEN_1950 & _GEN_1864;	// rob.scala:346:{27,69}, :347:31
    _GEN_1994 = _GEN_65 ? ~_GEN_1993 & _GEN_1866 : ~_GEN_1951 & _GEN_1866;	// rob.scala:346:{27,69}, :347:31
    _GEN_1996 = _GEN_65 ? ~_GEN_1995 & _GEN_1868 : ~_GEN_1952 & _GEN_1868;	// rob.scala:346:{27,69}, :347:31
    _GEN_1998 = _GEN_65 ? ~_GEN_1997 & _GEN_1870 : ~_GEN_1953 & _GEN_1870;	// rob.scala:346:{27,69}, :347:31
    _GEN_2000 = _GEN_65 ? ~_GEN_1999 & _GEN_1872 : ~_GEN_1954 & _GEN_1872;	// rob.scala:346:{27,69}, :347:31
    _GEN_2002 = _GEN_65 ? ~_GEN_2001 & _GEN_1874 : ~_GEN_1955 & _GEN_1874;	// rob.scala:346:{27,69}, :347:31
    _GEN_2004 = _GEN_65 ? ~_GEN_2003 & _GEN_1876 : ~_GEN_1956 & _GEN_1876;	// rob.scala:346:{27,69}, :347:31
    _GEN_2006 = _GEN_65 ? ~_GEN_2005 & _GEN_1878 : ~_GEN_1957 & _GEN_1878;	// rob.scala:346:{27,69}, :347:31
    _GEN_2008 = _GEN_65 ? ~_GEN_2007 & _GEN_1880 : ~_GEN_1958 & _GEN_1880;	// rob.scala:346:{27,69}, :347:31
    _GEN_2010 = _GEN_65 ? ~_GEN_2009 & _GEN_1882 : ~_GEN_1959 & _GEN_1882;	// rob.scala:346:{27,69}, :347:31
    _GEN_2012 = _GEN_65 ? ~_GEN_2011 & _GEN_1884 : ~_GEN_1960 & _GEN_1884;	// rob.scala:346:{27,69}, :347:31
    _GEN_2014 = _GEN_65 ? ~_GEN_2013 & _GEN_1886 : ~_GEN_1961 & _GEN_1886;	// rob.scala:346:{27,69}, :347:31
    _GEN_2016 = _GEN_65 ? ~_GEN_2015 & _GEN_1888 : ~_GEN_1962 & _GEN_1888;	// rob.scala:346:{27,69}, :347:31
    _GEN_2018 = _GEN_65 ? ~_GEN_2017 & _GEN_1890 : ~_GEN_1963 & _GEN_1890;	// rob.scala:346:{27,69}, :347:31
    _GEN_2020 = _GEN_65 ? ~_GEN_2019 & _GEN_1892 : ~_GEN_1964 & _GEN_1892;	// rob.scala:346:{27,69}, :347:31
    _GEN_2022 = _GEN_65 ? ~_GEN_2021 & _GEN_1894 : ~_GEN_1965 & _GEN_1894;	// rob.scala:346:{27,69}, :347:31
    _GEN_2024 = _GEN_65 ? ~_GEN_2023 & _GEN_1896 : ~_GEN_1966 & _GEN_1896;	// rob.scala:346:{27,69}, :347:31
    _GEN_2026 = _GEN_65 ? ~_GEN_2025 & _GEN_1898 : ~_GEN_1967 & _GEN_1898;	// rob.scala:346:{27,69}, :347:31
    _GEN_2028 = _GEN_65 ? ~_GEN_2027 & _GEN_1900 : ~_GEN_1968 & _GEN_1900;	// rob.scala:346:{27,69}, :347:31
    _GEN_2030 = _GEN_65 ? ~_GEN_2029 & _GEN_1902 : ~_GEN_1969 & _GEN_1902;	// rob.scala:346:{27,69}, :347:31
    _GEN_2032 = _GEN_65 ? ~_GEN_2031 & _GEN_1904 : ~_GEN_1970 & _GEN_1904;	// rob.scala:346:{27,69}, :347:31
    _GEN_2034 = _GEN_65 ? ~_GEN_2033 & _GEN_1906 : ~_GEN_1971 & _GEN_1906;	// rob.scala:346:{27,69}, :347:31
    _GEN_2036 = _GEN_65 ? ~_GEN_2035 & _GEN_1908 : ~_GEN_1972 & _GEN_1908;	// rob.scala:346:{27,69}, :347:31
    _GEN_2037 = _GEN_65 ? ~_GEN_1973 & _GEN_1909 : ~_GEN_1941 & _GEN_1909;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2038 = _GEN_65 ? ~_GEN_1975 & _GEN_1910 : ~_GEN_1942 & _GEN_1910;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2039 = _GEN_65 ? ~_GEN_1977 & _GEN_1911 : ~_GEN_1943 & _GEN_1911;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2040 = _GEN_65 ? ~_GEN_1979 & _GEN_1912 : ~_GEN_1944 & _GEN_1912;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2041 = _GEN_65 ? ~_GEN_1981 & _GEN_1913 : ~_GEN_1945 & _GEN_1913;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2042 = _GEN_65 ? ~_GEN_1983 & _GEN_1914 : ~_GEN_1946 & _GEN_1914;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2043 = _GEN_65 ? ~_GEN_1985 & _GEN_1915 : ~_GEN_1947 & _GEN_1915;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2044 = _GEN_65 ? ~_GEN_1987 & _GEN_1916 : ~_GEN_1948 & _GEN_1916;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2045 = _GEN_65 ? ~_GEN_1989 & _GEN_1917 : ~_GEN_1949 & _GEN_1917;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2046 = _GEN_65 ? ~_GEN_1991 & _GEN_1918 : ~_GEN_1950 & _GEN_1918;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2047 = _GEN_65 ? ~_GEN_1993 & _GEN_1919 : ~_GEN_1951 & _GEN_1919;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2048 = _GEN_65 ? ~_GEN_1995 & _GEN_1920 : ~_GEN_1952 & _GEN_1920;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2049 = _GEN_65 ? ~_GEN_1997 & _GEN_1921 : ~_GEN_1953 & _GEN_1921;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2050 = _GEN_65 ? ~_GEN_1999 & _GEN_1922 : ~_GEN_1954 & _GEN_1922;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2051 = _GEN_65 ? ~_GEN_2001 & _GEN_1923 : ~_GEN_1955 & _GEN_1923;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2052 = _GEN_65 ? ~_GEN_2003 & _GEN_1924 : ~_GEN_1956 & _GEN_1924;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2053 = _GEN_65 ? ~_GEN_2005 & _GEN_1925 : ~_GEN_1957 & _GEN_1925;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2054 = _GEN_65 ? ~_GEN_2007 & _GEN_1926 : ~_GEN_1958 & _GEN_1926;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2055 = _GEN_65 ? ~_GEN_2009 & _GEN_1927 : ~_GEN_1959 & _GEN_1927;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2056 = _GEN_65 ? ~_GEN_2011 & _GEN_1928 : ~_GEN_1960 & _GEN_1928;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2057 = _GEN_65 ? ~_GEN_2013 & _GEN_1929 : ~_GEN_1961 & _GEN_1929;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2058 = _GEN_65 ? ~_GEN_2015 & _GEN_1930 : ~_GEN_1962 & _GEN_1930;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2059 = _GEN_65 ? ~_GEN_2017 & _GEN_1931 : ~_GEN_1963 & _GEN_1931;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2060 = _GEN_65 ? ~_GEN_2019 & _GEN_1932 : ~_GEN_1964 & _GEN_1932;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2061 = _GEN_65 ? ~_GEN_2021 & _GEN_1933 : ~_GEN_1965 & _GEN_1933;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2062 = _GEN_65 ? ~_GEN_2023 & _GEN_1934 : ~_GEN_1966 & _GEN_1934;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2063 = _GEN_65 ? ~_GEN_2025 & _GEN_1935 : ~_GEN_1967 & _GEN_1935;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2064 = _GEN_65 ? ~_GEN_2027 & _GEN_1936 : ~_GEN_1968 & _GEN_1936;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2065 = _GEN_65 ? ~_GEN_2029 & _GEN_1937 : ~_GEN_1969 & _GEN_1937;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2066 = _GEN_65 ? ~_GEN_2031 & _GEN_1938 : ~_GEN_1970 & _GEN_1938;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2067 = _GEN_65 ? ~_GEN_2033 & _GEN_1939 : ~_GEN_1971 & _GEN_1939;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2068 = _GEN_65 ? ~_GEN_2035 & _GEN_1940 : ~_GEN_1972 & _GEN_1940;	// rob.scala:346:{27,69}, :347:31, :348:31
    _GEN_2069 = _GEN_66 & _GEN_793;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2070 = _GEN_66 & _GEN_795;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2071 = _GEN_66 & _GEN_797;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2072 = _GEN_66 & _GEN_799;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2073 = _GEN_66 & _GEN_801;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2074 = _GEN_66 & _GEN_803;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2075 = _GEN_66 & _GEN_805;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2076 = _GEN_66 & _GEN_807;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2077 = _GEN_66 & _GEN_809;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2078 = _GEN_66 & _GEN_811;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2079 = _GEN_66 & _GEN_813;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2080 = _GEN_66 & _GEN_815;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2081 = _GEN_66 & _GEN_817;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2082 = _GEN_66 & _GEN_819;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2083 = _GEN_66 & _GEN_821;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2084 = _GEN_66 & _GEN_823;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2085 = _GEN_66 & _GEN_825;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2086 = _GEN_66 & _GEN_827;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2087 = _GEN_66 & _GEN_829;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2088 = _GEN_66 & _GEN_831;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2089 = _GEN_66 & _GEN_833;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2090 = _GEN_66 & _GEN_835;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2091 = _GEN_66 & _GEN_837;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2092 = _GEN_66 & _GEN_839;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2093 = _GEN_66 & _GEN_841;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2094 = _GEN_66 & _GEN_843;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2095 = _GEN_66 & _GEN_845;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2096 = _GEN_66 & _GEN_847;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2097 = _GEN_66 & _GEN_849;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2098 = _GEN_66 & _GEN_851;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2099 = _GEN_66 & _GEN_853;	// rob.scala:346:69, :361:{31,75}, :363:26
    _GEN_2100 = _GEN_66 & (&(io_lsu_clr_bsy_0_bits[6:2]));	// rob.scala:236:31, :268:25, :346:69, :361:{31,75}, :363:26
    _GEN_2101 = rbk_row_2 & _GEN_918;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2102 = rbk_row_2 & _GEN_920;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2103 = rbk_row_2 & _GEN_922;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2104 = rbk_row_2 & _GEN_924;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2105 = rbk_row_2 & _GEN_926;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2106 = rbk_row_2 & _GEN_928;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2107 = rbk_row_2 & _GEN_930;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2108 = rbk_row_2 & _GEN_932;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2109 = rbk_row_2 & _GEN_934;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2110 = rbk_row_2 & _GEN_936;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2111 = rbk_row_2 & _GEN_938;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2112 = rbk_row_2 & _GEN_940;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2113 = rbk_row_2 & _GEN_942;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2114 = rbk_row_2 & _GEN_944;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2115 = rbk_row_2 & _GEN_946;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2116 = rbk_row_2 & _GEN_948;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2117 = rbk_row_2 & _GEN_950;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2118 = rbk_row_2 & _GEN_952;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2119 = rbk_row_2 & _GEN_954;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2120 = rbk_row_2 & _GEN_956;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2121 = rbk_row_2 & _GEN_958;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2122 = rbk_row_2 & _GEN_960;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2123 = rbk_row_2 & _GEN_962;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2124 = rbk_row_2 & _GEN_964;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2125 = rbk_row_2 & _GEN_966;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2126 = rbk_row_2 & _GEN_968;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2127 = rbk_row_2 & _GEN_970;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2128 = rbk_row_2 & _GEN_972;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2129 = rbk_row_2 & _GEN_974;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2130 = rbk_row_2 & _GEN_976;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2131 = rbk_row_2 & _GEN_978;	// rob.scala:323:29, :425:44, :433:20, :434:30
    _GEN_2132 = rbk_row_2 & (&com_idx);	// rob.scala:236:20, :323:29, :425:44, :433:20, :434:30
    _GEN_2133 = io_brupdate_b1_mispredict_mask & rob_uop_2_0_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2134 = io_brupdate_b1_mispredict_mask & rob_uop_2_1_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2135 = io_brupdate_b1_mispredict_mask & rob_uop_2_2_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2136 = io_brupdate_b1_mispredict_mask & rob_uop_2_3_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2137 = io_brupdate_b1_mispredict_mask & rob_uop_2_4_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2138 = io_brupdate_b1_mispredict_mask & rob_uop_2_5_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2139 = io_brupdate_b1_mispredict_mask & rob_uop_2_6_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2140 = io_brupdate_b1_mispredict_mask & rob_uop_2_7_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2141 = io_brupdate_b1_mispredict_mask & rob_uop_2_8_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2142 = io_brupdate_b1_mispredict_mask & rob_uop_2_9_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2143 = io_brupdate_b1_mispredict_mask & rob_uop_2_10_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2144 = io_brupdate_b1_mispredict_mask & rob_uop_2_11_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2145 = io_brupdate_b1_mispredict_mask & rob_uop_2_12_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2146 = io_brupdate_b1_mispredict_mask & rob_uop_2_13_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2147 = io_brupdate_b1_mispredict_mask & rob_uop_2_14_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2148 = io_brupdate_b1_mispredict_mask & rob_uop_2_15_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2149 = io_brupdate_b1_mispredict_mask & rob_uop_2_16_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2150 = io_brupdate_b1_mispredict_mask & rob_uop_2_17_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2151 = io_brupdate_b1_mispredict_mask & rob_uop_2_18_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2152 = io_brupdate_b1_mispredict_mask & rob_uop_2_19_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2153 = io_brupdate_b1_mispredict_mask & rob_uop_2_20_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2154 = io_brupdate_b1_mispredict_mask & rob_uop_2_21_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2155 = io_brupdate_b1_mispredict_mask & rob_uop_2_22_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2156 = io_brupdate_b1_mispredict_mask & rob_uop_2_23_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2157 = io_brupdate_b1_mispredict_mask & rob_uop_2_24_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2158 = io_brupdate_b1_mispredict_mask & rob_uop_2_25_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2159 = io_brupdate_b1_mispredict_mask & rob_uop_2_26_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2160 = io_brupdate_b1_mispredict_mask & rob_uop_2_27_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2161 = io_brupdate_b1_mispredict_mask & rob_uop_2_28_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2162 = io_brupdate_b1_mispredict_mask & rob_uop_2_29_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2163 = io_brupdate_b1_mispredict_mask & rob_uop_2_30_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2164 = io_brupdate_b1_mispredict_mask & rob_uop_2_31_br_mask;	// rob.scala:310:28, util.scala:118:51
    _GEN_2165 = ~(_io_flush_valid_output | exception_thrown) & rob_state != 2'h2;	// rob.scala:221:26, :236:31, :545:85, :573:36, :631:{9,26,47,60}
    _GEN_2166 =
      ~r_xcpt_val | io_lxcpt_bits_uop_rob_idx < r_xcpt_uop_rob_idx
      ^ io_lxcpt_bits_uop_rob_idx < rob_head_idx ^ r_xcpt_uop_rob_idx < rob_head_idx;	// Cat.scala:30:58, rob.scala:258:33, :259:29, :635:{13,25}, util.scala:363:{52,64,72,78}
    _GEN_2167 =
      ~r_xcpt_val
      & (enq_xcpts_0 | enq_xcpts_1 | io_enq_valids_2 & io_enq_uops_2_exception);	// rob.scala:258:33, :628:38, :635:13, :641:{30,51}
    idx = enq_xcpts_0 ? 2'h0 : enq_xcpts_1 ? 2'h1 : 2'h2;	// rob.scala:221:26, :236:31, :540:33, :628:38, :642:37
    next_xcpt_uop_br_mask =
      _GEN_2165
        ? (io_lxcpt_valid
             ? (_GEN_2166 ? io_lxcpt_bits_uop_br_mask : r_xcpt_uop_br_mask)
             : _GEN_2167 ? _GEN_2168[idx] : r_xcpt_uop_br_mask)
        : r_xcpt_uop_br_mask;	// rob.scala:259:29, :625:17, :631:{47,76}, :632:27, :635:{25,93}, :637:33, :641:{30,56}, :642:37, :646:23
    if (reset) begin
      rob_state <= 2'h0;	// rob.scala:221:26
      rob_head <= 5'h0;	// rob.scala:224:29
      rob_head_lsb <= 2'h0;	// rob.scala:221:26, :225:29
      rob_tail <= 5'h0;	// rob.scala:224:29, :228:29
      rob_tail_lsb <= 2'h0;	// rob.scala:221:26, :229:29
      rob_pnr <= 5'h0;	// rob.scala:224:29, :232:29
      rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
      maybe_full <= 1'h0;	// rob.scala:239:29, :361:75, :370:59, :372:26
      r_xcpt_val <= 1'h0;	// rob.scala:258:33, :361:75, :370:59, :372:26
      rob_val_0 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_3 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_4 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_5 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_6 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_7 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_8 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_9 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_10 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_11 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_12 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_13 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_14 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_15 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_16 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_17 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_18 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_19 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_20 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_21 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_22 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_23 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_24 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_25 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_26 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_27 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_28 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_29 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_30 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_31 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_0 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_1 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_2 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_3 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_4 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_5 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_6 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_7 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_8 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_9 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_10 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_11 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_12 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_13 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_14 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_15 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_16 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_17 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_18 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_19 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_20 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_21 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_22 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_23 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_24 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_25 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_26 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_27 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_28 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_29 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_30 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_1_31 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_0 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_1 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_2 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_3 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_4 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_5 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_6 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_7 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_8 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_9 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_10 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_11 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_12 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_13 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_14 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_15 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_16 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_17 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_18 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_19 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_20 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_21 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_22 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_23 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_24 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_25 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_26 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_27 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_28 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_29 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_30 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      rob_val_2_31 <= 1'h0;	// rob.scala:307:32, :361:75, :370:59, :372:26
      r_partial_row <= 1'h0;	// rob.scala:361:75, :370:59, :372:26, :677:30
      pnr_maybe_at_tail <= 1'h0;	// rob.scala:361:75, :370:59, :372:26, :714:36
    end
    else begin
      automatic logic            _GEN_2170;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2171;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2172;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2173;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2174;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2175;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2176;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2177;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2178;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2179;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2180;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2181;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2182;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2183;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2184;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2185;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2186;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2187;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2188;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2189;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2190;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2191;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2192;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2193;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2194;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2195;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2196;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2197;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2198;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2199;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2200;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2201;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2202;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2203;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2204;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2205;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2206;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2207;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2208;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2209;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2210;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2211;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2212;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2213;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2214;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2215;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2216;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2217;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2218;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2219;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2220;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2221;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2222;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2223;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2224;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2225;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2226;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2227;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2228;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2229;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2230;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2231;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2232;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2233;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2234;	// rob.scala:476:25
      automatic logic            _GEN_2235;	// rob.scala:476:25
      automatic logic            _GEN_2236;	// rob.scala:476:25
      automatic logic            _GEN_2237;	// rob.scala:476:25
      automatic logic            _GEN_2238;	// rob.scala:476:25
      automatic logic            _GEN_2239;	// rob.scala:476:25
      automatic logic            _GEN_2240;	// rob.scala:476:25
      automatic logic            _GEN_2241;	// rob.scala:476:25
      automatic logic            _GEN_2242;	// rob.scala:476:25
      automatic logic            _GEN_2243;	// rob.scala:476:25
      automatic logic            _GEN_2244;	// rob.scala:476:25
      automatic logic            _GEN_2245;	// rob.scala:476:25
      automatic logic            _GEN_2246;	// rob.scala:476:25
      automatic logic            _GEN_2247;	// rob.scala:476:25
      automatic logic            _GEN_2248;	// rob.scala:476:25
      automatic logic            _GEN_2249;	// rob.scala:476:25
      automatic logic            _GEN_2250;	// rob.scala:476:25
      automatic logic            _GEN_2251;	// rob.scala:476:25
      automatic logic            _GEN_2252;	// rob.scala:476:25
      automatic logic            _GEN_2253;	// rob.scala:476:25
      automatic logic            _GEN_2254;	// rob.scala:476:25
      automatic logic            _GEN_2255;	// rob.scala:476:25
      automatic logic            _GEN_2256;	// rob.scala:476:25
      automatic logic            _GEN_2257;	// rob.scala:476:25
      automatic logic            _GEN_2258;	// rob.scala:476:25
      automatic logic            _GEN_2259;	// rob.scala:476:25
      automatic logic            _GEN_2260;	// rob.scala:476:25
      automatic logic            _GEN_2261;	// rob.scala:476:25
      automatic logic            _GEN_2262;	// rob.scala:476:25
      automatic logic            _GEN_2263;	// rob.scala:476:25
      automatic logic            _GEN_2264;	// rob.scala:476:25
      automatic logic            rob_pnr_unsafe_0;	// rob.scala:493:43
      automatic logic            _GEN_2265;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2266;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2267;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2268;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2269;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2270;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2271;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2272;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2273;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2274;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2275;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2276;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2277;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2278;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2279;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2280;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2281;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2282;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2283;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2284;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2285;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2286;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2287;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2288;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2289;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2290;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2291;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2292;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2293;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2294;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2295;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2296;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2297;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2298;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2299;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2300;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2301;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2302;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2303;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2304;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2305;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2306;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2307;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2308;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2309;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2310;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2311;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2312;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2313;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2314;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2315;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2316;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2317;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2318;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2319;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2320;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2321;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2322;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2323;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2324;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2325;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2326;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2327;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2328;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            rob_pnr_unsafe_1;	// rob.scala:493:43
      automatic logic            _GEN_2329;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2330;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2331;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2332;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2333;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2334;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2335;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2336;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2337;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2338;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2339;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2340;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2341;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2342;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2343;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2344;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2345;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2346;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2347;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2348;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2349;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2350;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2351;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2352;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2353;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2354;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2355;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2356;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2357;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2358;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2359;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2360;	// rob.scala:307:32, :323:29, :324:31
      automatic logic            _GEN_2361;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2362;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2363;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2364;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2365;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2366;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2367;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2368;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2369;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2370;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2371;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2372;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2373;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2374;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2375;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2376;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2377;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2378;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2379;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2380;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2381;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2382;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2383;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2384;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2385;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2386;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2387;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2388;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2389;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2390;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2391;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _GEN_2392;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20
      automatic logic            _do_inc_row_T_3;	// rob.scala:717:64
      automatic logic            do_inc_row;	// rob.scala:717:52
      automatic logic [2:0]      _GEN_2393;	// rob.scala:718:34
      automatic logic            _GEN_2394;	// rob.scala:755:68
      automatic logic            _GEN_2395;	// rob.scala:761:45
      automatic logic [1:0]      _GEN_2396;	// rob.scala:221:26, :819:22, :820:21
      automatic logic [3:0][1:0] _GEN_2397;	// Conditional.scala:37:30, :39:67, :40:58, rob.scala:221:26, :540:61, :804:19, :808:51, :819:22, :824:42
      _GEN_2170 = _GEN_97 | rob_val_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2171 = _GEN_99 | rob_val_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2172 = _GEN_101 | rob_val_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2173 = _GEN_103 | rob_val_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2174 = _GEN_105 | rob_val_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2175 = _GEN_107 | rob_val_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2176 = _GEN_109 | rob_val_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2177 = _GEN_111 | rob_val_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2178 = _GEN_113 | rob_val_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2179 = _GEN_115 | rob_val_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2180 = _GEN_117 | rob_val_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2181 = _GEN_119 | rob_val_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2182 = _GEN_121 | rob_val_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2183 = _GEN_123 | rob_val_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2184 = _GEN_125 | rob_val_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2185 = _GEN_127 | rob_val_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2186 = _GEN_129 | rob_val_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2187 = _GEN_131 | rob_val_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2188 = _GEN_133 | rob_val_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2189 = _GEN_135 | rob_val_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2190 = _GEN_137 | rob_val_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2191 = _GEN_139 | rob_val_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2192 = _GEN_141 | rob_val_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2193 = _GEN_143 | rob_val_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2194 = _GEN_145 | rob_val_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2195 = _GEN_147 | rob_val_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2196 = _GEN_149 | rob_val_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2197 = _GEN_151 | rob_val_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2198 = _GEN_153 | rob_val_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2199 = _GEN_155 | rob_val_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2200 = _GEN_157 | rob_val_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2201 = _GEN_158 | rob_val_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2202 = (|_GEN_981) | _GEN_919;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2203 = (|_GEN_982) | _GEN_921;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2204 = (|_GEN_983) | _GEN_923;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2205 = (|_GEN_984) | _GEN_925;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2206 = (|_GEN_985) | _GEN_927;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2207 = (|_GEN_986) | _GEN_929;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2208 = (|_GEN_987) | _GEN_931;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2209 = (|_GEN_988) | _GEN_933;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2210 = (|_GEN_989) | _GEN_935;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2211 = (|_GEN_990) | _GEN_937;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2212 = (|_GEN_991) | _GEN_939;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2213 = (|_GEN_992) | _GEN_941;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2214 = (|_GEN_993) | _GEN_943;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2215 = (|_GEN_994) | _GEN_945;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2216 = (|_GEN_995) | _GEN_947;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2217 = (|_GEN_996) | _GEN_949;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2218 = (|_GEN_997) | _GEN_951;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2219 = (|_GEN_998) | _GEN_953;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2220 = (|_GEN_999) | _GEN_955;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2221 = (|_GEN_1000) | _GEN_957;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2222 = (|_GEN_1001) | _GEN_959;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2223 = (|_GEN_1002) | _GEN_961;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2224 = (|_GEN_1003) | _GEN_963;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2225 = (|_GEN_1004) | _GEN_965;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2226 = (|_GEN_1005) | _GEN_967;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2227 = (|_GEN_1006) | _GEN_969;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2228 = (|_GEN_1007) | _GEN_971;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2229 = (|_GEN_1008) | _GEN_973;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2230 = (|_GEN_1009) | _GEN_975;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2231 = (|_GEN_1010) | _GEN_977;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2232 = (|_GEN_1011) | _GEN_979;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2233 = (|_GEN_1012) | _GEN_980;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2234 = rob_head == 5'h0;	// rob.scala:224:29, :476:25
      _GEN_2235 = rob_head == 5'h1;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2236 = rob_head == 5'h2;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2237 = rob_head == 5'h3;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2238 = rob_head == 5'h4;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2239 = rob_head == 5'h5;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2240 = rob_head == 5'h6;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2241 = rob_head == 5'h7;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2242 = rob_head == 5'h8;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2243 = rob_head == 5'h9;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2244 = rob_head == 5'hA;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2245 = rob_head == 5'hB;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2246 = rob_head == 5'hC;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2247 = rob_head == 5'hD;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2248 = rob_head == 5'hE;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2249 = rob_head == 5'hF;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2250 = rob_head == 5'h10;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2251 = rob_head == 5'h11;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2252 = rob_head == 5'h12;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2253 = rob_head == 5'h13;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2254 = rob_head == 5'h14;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2255 = rob_head == 5'h15;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2256 = rob_head == 5'h16;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2257 = rob_head == 5'h17;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2258 = rob_head == 5'h18;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2259 = rob_head == 5'h19;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2260 = rob_head == 5'h1A;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2261 = rob_head == 5'h1B;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2262 = rob_head == 5'h1C;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2263 = rob_head == 5'h1D;	// rob.scala:224:29, :324:31, :476:25
      _GEN_2264 = rob_head == 5'h1E;	// rob.scala:224:29, :324:31, :476:25
      rob_pnr_unsafe_0 = _GEN[rob_pnr] & (_GEN_10[rob_pnr] | _GEN_11[rob_pnr]);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}
      _GEN_2265 = _GEN_1013 | rob_val_1_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2266 = _GEN_1014 | rob_val_1_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2267 = _GEN_1015 | rob_val_1_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2268 = _GEN_1016 | rob_val_1_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2269 = _GEN_1017 | rob_val_1_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2270 = _GEN_1018 | rob_val_1_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2271 = _GEN_1019 | rob_val_1_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2272 = _GEN_1020 | rob_val_1_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2273 = _GEN_1021 | rob_val_1_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2274 = _GEN_1022 | rob_val_1_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2275 = _GEN_1023 | rob_val_1_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2276 = _GEN_1024 | rob_val_1_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2277 = _GEN_1025 | rob_val_1_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2278 = _GEN_1026 | rob_val_1_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2279 = _GEN_1027 | rob_val_1_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2280 = _GEN_1028 | rob_val_1_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2281 = _GEN_1029 | rob_val_1_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2282 = _GEN_1030 | rob_val_1_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2283 = _GEN_1031 | rob_val_1_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2284 = _GEN_1032 | rob_val_1_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2285 = _GEN_1033 | rob_val_1_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2286 = _GEN_1034 | rob_val_1_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2287 = _GEN_1035 | rob_val_1_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2288 = _GEN_1036 | rob_val_1_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2289 = _GEN_1037 | rob_val_1_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2290 = _GEN_1038 | rob_val_1_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2291 = _GEN_1039 | rob_val_1_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2292 = _GEN_1040 | rob_val_1_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2293 = _GEN_1041 | rob_val_1_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2294 = _GEN_1042 | rob_val_1_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2295 = _GEN_1043 | rob_val_1_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2296 = _GEN_1044 | rob_val_1_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2297 = (|_GEN_1557) | _GEN_1525;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2298 = (|_GEN_1558) | _GEN_1526;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2299 = (|_GEN_1559) | _GEN_1527;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2300 = (|_GEN_1560) | _GEN_1528;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2301 = (|_GEN_1561) | _GEN_1529;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2302 = (|_GEN_1562) | _GEN_1530;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2303 = (|_GEN_1563) | _GEN_1531;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2304 = (|_GEN_1564) | _GEN_1532;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2305 = (|_GEN_1565) | _GEN_1533;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2306 = (|_GEN_1566) | _GEN_1534;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2307 = (|_GEN_1567) | _GEN_1535;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2308 = (|_GEN_1568) | _GEN_1536;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2309 = (|_GEN_1569) | _GEN_1537;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2310 = (|_GEN_1570) | _GEN_1538;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2311 = (|_GEN_1571) | _GEN_1539;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2312 = (|_GEN_1572) | _GEN_1540;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2313 = (|_GEN_1573) | _GEN_1541;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2314 = (|_GEN_1574) | _GEN_1542;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2315 = (|_GEN_1575) | _GEN_1543;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2316 = (|_GEN_1576) | _GEN_1544;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2317 = (|_GEN_1577) | _GEN_1545;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2318 = (|_GEN_1578) | _GEN_1546;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2319 = (|_GEN_1579) | _GEN_1547;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2320 = (|_GEN_1580) | _GEN_1548;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2321 = (|_GEN_1581) | _GEN_1549;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2322 = (|_GEN_1582) | _GEN_1550;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2323 = (|_GEN_1583) | _GEN_1551;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2324 = (|_GEN_1584) | _GEN_1552;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2325 = (|_GEN_1585) | _GEN_1553;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2326 = (|_GEN_1586) | _GEN_1554;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2327 = (|_GEN_1587) | _GEN_1555;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2328 = (|_GEN_1588) | _GEN_1556;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      rob_pnr_unsafe_1 = _GEN_29[rob_pnr] & (_GEN_40[rob_pnr] | _GEN_41[rob_pnr]);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}
      _GEN_2329 = _GEN_1589 | rob_val_2_0;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2330 = _GEN_1590 | rob_val_2_1;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2331 = _GEN_1591 | rob_val_2_2;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2332 = _GEN_1592 | rob_val_2_3;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2333 = _GEN_1593 | rob_val_2_4;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2334 = _GEN_1594 | rob_val_2_5;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2335 = _GEN_1595 | rob_val_2_6;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2336 = _GEN_1596 | rob_val_2_7;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2337 = _GEN_1597 | rob_val_2_8;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2338 = _GEN_1598 | rob_val_2_9;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2339 = _GEN_1599 | rob_val_2_10;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2340 = _GEN_1600 | rob_val_2_11;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2341 = _GEN_1601 | rob_val_2_12;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2342 = _GEN_1602 | rob_val_2_13;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2343 = _GEN_1603 | rob_val_2_14;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2344 = _GEN_1604 | rob_val_2_15;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2345 = _GEN_1605 | rob_val_2_16;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2346 = _GEN_1606 | rob_val_2_17;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2347 = _GEN_1607 | rob_val_2_18;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2348 = _GEN_1608 | rob_val_2_19;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2349 = _GEN_1609 | rob_val_2_20;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2350 = _GEN_1610 | rob_val_2_21;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2351 = _GEN_1611 | rob_val_2_22;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2352 = _GEN_1612 | rob_val_2_23;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2353 = _GEN_1613 | rob_val_2_24;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2354 = _GEN_1614 | rob_val_2_25;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2355 = _GEN_1615 | rob_val_2_26;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2356 = _GEN_1616 | rob_val_2_27;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2357 = _GEN_1617 | rob_val_2_28;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2358 = _GEN_1618 | rob_val_2_29;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2359 = _GEN_1619 | rob_val_2_30;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2360 = _GEN_1620 | rob_val_2_31;	// rob.scala:307:32, :323:29, :324:31
      _GEN_2361 = (|_GEN_2133) | _GEN_2101;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2362 = (|_GEN_2134) | _GEN_2102;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2363 = (|_GEN_2135) | _GEN_2103;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2364 = (|_GEN_2136) | _GEN_2104;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2365 = (|_GEN_2137) | _GEN_2105;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2366 = (|_GEN_2138) | _GEN_2106;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2367 = (|_GEN_2139) | _GEN_2107;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2368 = (|_GEN_2140) | _GEN_2108;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2369 = (|_GEN_2141) | _GEN_2109;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2370 = (|_GEN_2142) | _GEN_2110;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2371 = (|_GEN_2143) | _GEN_2111;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2372 = (|_GEN_2144) | _GEN_2112;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2373 = (|_GEN_2145) | _GEN_2113;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2374 = (|_GEN_2146) | _GEN_2114;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2375 = (|_GEN_2147) | _GEN_2115;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2376 = (|_GEN_2148) | _GEN_2116;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2377 = (|_GEN_2149) | _GEN_2117;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2378 = (|_GEN_2150) | _GEN_2118;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2379 = (|_GEN_2151) | _GEN_2119;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2380 = (|_GEN_2152) | _GEN_2120;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2381 = (|_GEN_2153) | _GEN_2121;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2382 = (|_GEN_2154) | _GEN_2122;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2383 = (|_GEN_2155) | _GEN_2123;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2384 = (|_GEN_2156) | _GEN_2124;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2385 = (|_GEN_2157) | _GEN_2125;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2386 = (|_GEN_2158) | _GEN_2126;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2387 = (|_GEN_2159) | _GEN_2127;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2388 = (|_GEN_2160) | _GEN_2128;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2389 = (|_GEN_2161) | _GEN_2129;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2390 = (|_GEN_2162) | _GEN_2130;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2391 = (|_GEN_2163) | _GEN_2131;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _GEN_2392 = (|_GEN_2164) | _GEN_2132;	// rob.scala:323:29, :433:20, :434:30, :455:7, :456:20, util.scala:118:{51,59}
      _do_inc_row_T_3 = rob_pnr != rob_tail;	// rob.scala:228:29, :232:29, :717:64
      do_inc_row =
        ~(rob_pnr_unsafe_0 | rob_pnr_unsafe_1 | _GEN_59[rob_pnr]
          & (_GEN_70[rob_pnr] | _GEN_71[rob_pnr]))
        & (_do_inc_row_T_3 | full & ~pnr_maybe_at_tail);	// rob.scala:232:29, :324:31, :394:15, :398:49, :493:{43,67}, :714:36, :717:{23,47,52,64,77,86,89}, :787:39
      _GEN_2393 = {io_enq_valids_2, io_enq_valids_1, io_enq_valids_0};	// rob.scala:718:34
      _GEN_2394 = _io_commit_rollback_T_2 & rob_tail == rob_head & ~maybe_full;	// rob.scala:224:29, :228:29, :236:31, :239:29, :686:49, :755:{54,68}
      _GEN_2395 = (|_GEN_2393) & ~io_enq_partial_stall;	// rob.scala:718:{34,41}, :761:{45,48}
      _GEN_2396 = empty ? 2'h1 : rob_state;	// rob.scala:221:26, :540:33, :788:41, :819:22, :820:21
      _GEN_2397 =
        {{REG_2 ? 2'h2 : _GEN_2396},
         {_GEN_2396},
         {REG_1
            ? 2'h2
            : io_enq_valids_2 & io_enq_uops_2_is_unique | io_enq_valids_1
              & io_enq_uops_1_is_unique | io_enq_valids_0 & io_enq_uops_0_is_unique
                ? 2'h3
                : rob_state},
         {2'h1}};	// Conditional.scala:37:30, :39:67, :40:58, rob.scala:221:26, :236:31, :419:36, :540:{33,61}, :804:19, :808:{22,51}, :809:21, :812:{36,65}, :813:25, :819:22, :820:21, :824:{22,42}, :825:21, :826:29
      rob_state <= _GEN_2397[rob_state];	// Conditional.scala:37:30, :39:67, :40:58, rob.scala:221:26, :540:61, :804:19, :808:51, :819:22, :824:42
      if (finished_committing_row)	// rob.scala:685:59
        rob_head <= rob_head + 5'h1;	// rob.scala:224:29, :324:31, util.scala:203:14
      if (finished_committing_row | rob_head_vals_0)	// rob.scala:398:49, :685:59, :688:34, :690:18, :693:18
        rob_head_lsb <= 2'h0;	// rob.scala:221:26, :225:29
      else	// rob.scala:688:34, :690:18, :693:18
        rob_head_lsb <= rob_head_vals_1 ? 2'h1 : {rob_head_vals_2, 1'h0};	// Mux.scala:47:69, rob.scala:225:29, :361:75, :370:59, :372:26, :398:49, :540:33
      if (_GEN_95) begin	// rob.scala:750:34
        rob_tail <= rob_tail - 5'h1;	// rob.scala:228:29, util.scala:220:14
        rob_tail_lsb <= 2'h2;	// rob.scala:229:29, :236:31
      end
      else if (_GEN_2394)	// rob.scala:755:68
        rob_tail_lsb <= rob_head_lsb;	// rob.scala:225:29, :229:29
      else begin	// rob.scala:755:68
        if (io_brupdate_b2_mispredict)
          rob_tail <= io_brupdate_b2_uop_rob_idx[6:2] + 5'h1;	// rob.scala:228:29, :236:31, :268:25, :324:31, util.scala:203:14
        else if (_GEN_2395)	// rob.scala:761:45
          rob_tail <= rob_tail + 5'h1;	// rob.scala:228:29, :324:31, util.scala:203:14
        if (io_brupdate_b2_mispredict | _GEN_2395)	// rob.scala:758:43, :760:18, :761:{45,71}, :763:18, :765:70
          rob_tail_lsb <= 2'h0;	// rob.scala:221:26, :229:29
        else if ((|_GEN_2393) & io_enq_partial_stall) begin	// rob.scala:718:{34,41}, :765:45
          automatic logic [1:0] _GEN_2398 =
            {io_enq_valids_1, io_enq_valids_0} | {io_enq_valids_2, io_enq_valids_1};	// util.scala:373:{29,45}
          automatic logic [1:0] _lo_T_37;	// rob.scala:766:37
          _lo_T_37 = ~{_GEN_2398[1], _GEN_2398[0] | io_enq_valids_2};	// rob.scala:236:31, :766:37, util.scala:373:{29,45}
          if (_lo_T_37[0])	// OneHot.scala:47:40, rob.scala:766:37
            rob_tail_lsb <= 2'h0;	// rob.scala:221:26, :229:29
          else if (_lo_T_37[1])	// OneHot.scala:47:40, rob.scala:766:37
            rob_tail_lsb <= 2'h1;	// rob.scala:229:29, :540:33
          else	// OneHot.scala:47:40
            rob_tail_lsb <= 2'h2;	// rob.scala:229:29, :236:31
        end
      end
      if (empty & (|_GEN_2393)) begin	// rob.scala:718:{17,34,41}, :788:41
        rob_pnr <= rob_head;	// rob.scala:224:29, :232:29
        if (io_enq_valids_0)
          rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
        else if (io_enq_valids_1)
          rob_pnr_lsb <= 2'h1;	// rob.scala:233:29, :540:33
        else
          rob_pnr_lsb <= 2'h2;	// rob.scala:233:29, :236:31
      end
      else begin	// rob.scala:718:17
        automatic logic safe_to_inc;	// rob.scala:716:46
        safe_to_inc = _io_ready_T | (&rob_state);	// rob.scala:221:26, :716:{33,46,59}
        if (safe_to_inc & do_inc_row) begin	// rob.scala:716:46, :717:52, :725:30
          rob_pnr <= rob_pnr + 5'h1;	// rob.scala:232:29, :324:31, util.scala:203:14
          rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
        end
        else if (safe_to_inc & (_do_inc_row_T_3 | full & ~pnr_maybe_at_tail)) begin	// rob.scala:714:36, :716:46, :717:{64,89}, :728:{30,55,64}, :787:39
          if (rob_pnr_unsafe_0)	// rob.scala:493:43
            rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
          else if (rob_pnr_unsafe_1)	// rob.scala:493:43
            rob_pnr_lsb <= 2'h1;	// rob.scala:233:29, :540:33
          else	// rob.scala:493:43
            rob_pnr_lsb <= 2'h2;	// rob.scala:233:29, :236:31
        end
        else if (safe_to_inc & ~full & ~empty) begin	// rob.scala:425:47, :716:46, :730:{39,42}, :787:39, :788:41
          automatic logic [1:0] _GEN_2399 =
            {rob_tail_vals_1, rob_tail_vals_0} | {rob_tail_vals_2, rob_tail_vals_1};	// rob.scala:324:31, util.scala:373:{29,45}
          automatic logic [1:0] _lo_T_25;	// rob.scala:731:60
          _lo_T_25 =
            {rob_pnr_unsafe_1, rob_pnr_unsafe_0}
            | ~{_GEN_2399[1], _GEN_2399[0] | rob_tail_vals_2};	// rob.scala:236:31, :324:31, :493:43, :731:{53,60,62}, util.scala:373:{29,45}
          if (_lo_T_25[0])	// OneHot.scala:47:40, rob.scala:731:60
            rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
          else if (_lo_T_25[1])	// OneHot.scala:47:40, rob.scala:731:60
            rob_pnr_lsb <= 2'h1;	// rob.scala:233:29, :540:33
          else	// OneHot.scala:47:40
            rob_pnr_lsb <= 2'h2;	// rob.scala:233:29, :236:31
        end
        else if (full & pnr_maybe_at_tail)	// rob.scala:714:36, :732:23, :787:39
          rob_pnr_lsb <= 2'h0;	// rob.scala:221:26, :233:29
      end
      maybe_full <=
        ~rob_deq
        & (~(_GEN_95 | _GEN_2394 | io_brupdate_b2_mispredict) & _GEN_2395 | maybe_full)
        | (|io_brupdate_b1_mispredict_mask);	// rob.scala:239:29, :688:34, :736:26, :750:{34,76}, :754:13, :755:{68,84}, :758:43, :761:{45,71}, :786:{26,38,53,87}
      r_xcpt_val <=
        ~(_io_flush_valid_output
          | (|(io_brupdate_b1_mispredict_mask & next_xcpt_uop_br_mask)))
        & (_GEN_2165
             ? (io_lxcpt_valid ? _GEN_2166 | r_xcpt_val : _GEN_2167 | r_xcpt_val)
             : r_xcpt_val);	// rob.scala:258:33, :573:36, :625:17, :631:{47,76}, :632:27, :635:{25,93}, :636:33, :641:{30,56}, :645:23, :654:{24,73}, :655:16, util.scala:118:{51,59}
      if (will_commit_0) begin	// rob.scala:547:70
        rob_val_0 <= ~(_GEN_2234 | _GEN_2202) & _GEN_2170;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1 <= ~(_GEN_2235 | _GEN_2203) & _GEN_2171;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2 <= ~(_GEN_2236 | _GEN_2204) & _GEN_2172;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_3 <= ~(_GEN_2237 | _GEN_2205) & _GEN_2173;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_4 <= ~(_GEN_2238 | _GEN_2206) & _GEN_2174;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_5 <= ~(_GEN_2239 | _GEN_2207) & _GEN_2175;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_6 <= ~(_GEN_2240 | _GEN_2208) & _GEN_2176;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_7 <= ~(_GEN_2241 | _GEN_2209) & _GEN_2177;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_8 <= ~(_GEN_2242 | _GEN_2210) & _GEN_2178;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_9 <= ~(_GEN_2243 | _GEN_2211) & _GEN_2179;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_10 <= ~(_GEN_2244 | _GEN_2212) & _GEN_2180;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_11 <= ~(_GEN_2245 | _GEN_2213) & _GEN_2181;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_12 <= ~(_GEN_2246 | _GEN_2214) & _GEN_2182;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_13 <= ~(_GEN_2247 | _GEN_2215) & _GEN_2183;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_14 <= ~(_GEN_2248 | _GEN_2216) & _GEN_2184;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_15 <= ~(_GEN_2249 | _GEN_2217) & _GEN_2185;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_16 <= ~(_GEN_2250 | _GEN_2218) & _GEN_2186;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_17 <= ~(_GEN_2251 | _GEN_2219) & _GEN_2187;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_18 <= ~(_GEN_2252 | _GEN_2220) & _GEN_2188;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_19 <= ~(_GEN_2253 | _GEN_2221) & _GEN_2189;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_20 <= ~(_GEN_2254 | _GEN_2222) & _GEN_2190;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_21 <= ~(_GEN_2255 | _GEN_2223) & _GEN_2191;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_22 <= ~(_GEN_2256 | _GEN_2224) & _GEN_2192;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_23 <= ~(_GEN_2257 | _GEN_2225) & _GEN_2193;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_24 <= ~(_GEN_2258 | _GEN_2226) & _GEN_2194;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_25 <= ~(_GEN_2259 | _GEN_2227) & _GEN_2195;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_26 <= ~(_GEN_2260 | _GEN_2228) & _GEN_2196;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_27 <= ~(_GEN_2261 | _GEN_2229) & _GEN_2197;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_28 <= ~(_GEN_2262 | _GEN_2230) & _GEN_2198;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_29 <= ~(_GEN_2263 | _GEN_2231) & _GEN_2199;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_30 <= ~(_GEN_2264 | _GEN_2232) & _GEN_2200;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_31 <= ~((&rob_head) | _GEN_2233) & _GEN_2201;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_0 <= ~_GEN_2202 & _GEN_2170;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1 <= ~_GEN_2203 & _GEN_2171;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2 <= ~_GEN_2204 & _GEN_2172;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_3 <= ~_GEN_2205 & _GEN_2173;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_4 <= ~_GEN_2206 & _GEN_2174;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_5 <= ~_GEN_2207 & _GEN_2175;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_6 <= ~_GEN_2208 & _GEN_2176;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_7 <= ~_GEN_2209 & _GEN_2177;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_8 <= ~_GEN_2210 & _GEN_2178;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_9 <= ~_GEN_2211 & _GEN_2179;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_10 <= ~_GEN_2212 & _GEN_2180;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_11 <= ~_GEN_2213 & _GEN_2181;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_12 <= ~_GEN_2214 & _GEN_2182;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_13 <= ~_GEN_2215 & _GEN_2183;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_14 <= ~_GEN_2216 & _GEN_2184;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_15 <= ~_GEN_2217 & _GEN_2185;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_16 <= ~_GEN_2218 & _GEN_2186;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_17 <= ~_GEN_2219 & _GEN_2187;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_18 <= ~_GEN_2220 & _GEN_2188;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_19 <= ~_GEN_2221 & _GEN_2189;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_20 <= ~_GEN_2222 & _GEN_2190;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_21 <= ~_GEN_2223 & _GEN_2191;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_22 <= ~_GEN_2224 & _GEN_2192;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_23 <= ~_GEN_2225 & _GEN_2193;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_24 <= ~_GEN_2226 & _GEN_2194;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_25 <= ~_GEN_2227 & _GEN_2195;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_26 <= ~_GEN_2228 & _GEN_2196;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_27 <= ~_GEN_2229 & _GEN_2197;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_28 <= ~_GEN_2230 & _GEN_2198;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_29 <= ~_GEN_2231 & _GEN_2199;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_30 <= ~_GEN_2232 & _GEN_2200;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_31 <= ~_GEN_2233 & _GEN_2201;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (will_commit_1) begin	// rob.scala:547:70
        rob_val_1_0 <= ~(_GEN_2234 | _GEN_2297) & _GEN_2265;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_1 <= ~(_GEN_2235 | _GEN_2298) & _GEN_2266;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_2 <= ~(_GEN_2236 | _GEN_2299) & _GEN_2267;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_3 <= ~(_GEN_2237 | _GEN_2300) & _GEN_2268;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_4 <= ~(_GEN_2238 | _GEN_2301) & _GEN_2269;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_5 <= ~(_GEN_2239 | _GEN_2302) & _GEN_2270;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_6 <= ~(_GEN_2240 | _GEN_2303) & _GEN_2271;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_7 <= ~(_GEN_2241 | _GEN_2304) & _GEN_2272;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_8 <= ~(_GEN_2242 | _GEN_2305) & _GEN_2273;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_9 <= ~(_GEN_2243 | _GEN_2306) & _GEN_2274;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_10 <= ~(_GEN_2244 | _GEN_2307) & _GEN_2275;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_11 <= ~(_GEN_2245 | _GEN_2308) & _GEN_2276;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_12 <= ~(_GEN_2246 | _GEN_2309) & _GEN_2277;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_13 <= ~(_GEN_2247 | _GEN_2310) & _GEN_2278;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_14 <= ~(_GEN_2248 | _GEN_2311) & _GEN_2279;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_15 <= ~(_GEN_2249 | _GEN_2312) & _GEN_2280;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_16 <= ~(_GEN_2250 | _GEN_2313) & _GEN_2281;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_17 <= ~(_GEN_2251 | _GEN_2314) & _GEN_2282;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_18 <= ~(_GEN_2252 | _GEN_2315) & _GEN_2283;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_19 <= ~(_GEN_2253 | _GEN_2316) & _GEN_2284;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_20 <= ~(_GEN_2254 | _GEN_2317) & _GEN_2285;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_21 <= ~(_GEN_2255 | _GEN_2318) & _GEN_2286;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_22 <= ~(_GEN_2256 | _GEN_2319) & _GEN_2287;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_23 <= ~(_GEN_2257 | _GEN_2320) & _GEN_2288;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_24 <= ~(_GEN_2258 | _GEN_2321) & _GEN_2289;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_25 <= ~(_GEN_2259 | _GEN_2322) & _GEN_2290;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_26 <= ~(_GEN_2260 | _GEN_2323) & _GEN_2291;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_27 <= ~(_GEN_2261 | _GEN_2324) & _GEN_2292;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_28 <= ~(_GEN_2262 | _GEN_2325) & _GEN_2293;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_29 <= ~(_GEN_2263 | _GEN_2326) & _GEN_2294;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_30 <= ~(_GEN_2264 | _GEN_2327) & _GEN_2295;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_1_31 <= ~((&rob_head) | _GEN_2328) & _GEN_2296;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_1_0 <= ~_GEN_2297 & _GEN_2265;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_1 <= ~_GEN_2298 & _GEN_2266;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_2 <= ~_GEN_2299 & _GEN_2267;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_3 <= ~_GEN_2300 & _GEN_2268;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_4 <= ~_GEN_2301 & _GEN_2269;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_5 <= ~_GEN_2302 & _GEN_2270;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_6 <= ~_GEN_2303 & _GEN_2271;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_7 <= ~_GEN_2304 & _GEN_2272;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_8 <= ~_GEN_2305 & _GEN_2273;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_9 <= ~_GEN_2306 & _GEN_2274;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_10 <= ~_GEN_2307 & _GEN_2275;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_11 <= ~_GEN_2308 & _GEN_2276;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_12 <= ~_GEN_2309 & _GEN_2277;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_13 <= ~_GEN_2310 & _GEN_2278;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_14 <= ~_GEN_2311 & _GEN_2279;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_15 <= ~_GEN_2312 & _GEN_2280;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_16 <= ~_GEN_2313 & _GEN_2281;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_17 <= ~_GEN_2314 & _GEN_2282;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_18 <= ~_GEN_2315 & _GEN_2283;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_19 <= ~_GEN_2316 & _GEN_2284;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_20 <= ~_GEN_2317 & _GEN_2285;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_21 <= ~_GEN_2318 & _GEN_2286;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_22 <= ~_GEN_2319 & _GEN_2287;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_23 <= ~_GEN_2320 & _GEN_2288;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_24 <= ~_GEN_2321 & _GEN_2289;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_25 <= ~_GEN_2322 & _GEN_2290;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_26 <= ~_GEN_2323 & _GEN_2291;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_27 <= ~_GEN_2324 & _GEN_2292;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_28 <= ~_GEN_2325 & _GEN_2293;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_29 <= ~_GEN_2326 & _GEN_2294;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_30 <= ~_GEN_2327 & _GEN_2295;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_1_31 <= ~_GEN_2328 & _GEN_2296;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (will_commit_2) begin	// rob.scala:547:70
        rob_val_2_0 <= ~(_GEN_2234 | _GEN_2361) & _GEN_2329;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_1 <= ~(_GEN_2235 | _GEN_2362) & _GEN_2330;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_2 <= ~(_GEN_2236 | _GEN_2363) & _GEN_2331;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_3 <= ~(_GEN_2237 | _GEN_2364) & _GEN_2332;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_4 <= ~(_GEN_2238 | _GEN_2365) & _GEN_2333;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_5 <= ~(_GEN_2239 | _GEN_2366) & _GEN_2334;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_6 <= ~(_GEN_2240 | _GEN_2367) & _GEN_2335;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_7 <= ~(_GEN_2241 | _GEN_2368) & _GEN_2336;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_8 <= ~(_GEN_2242 | _GEN_2369) & _GEN_2337;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_9 <= ~(_GEN_2243 | _GEN_2370) & _GEN_2338;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_10 <= ~(_GEN_2244 | _GEN_2371) & _GEN_2339;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_11 <= ~(_GEN_2245 | _GEN_2372) & _GEN_2340;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_12 <= ~(_GEN_2246 | _GEN_2373) & _GEN_2341;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_13 <= ~(_GEN_2247 | _GEN_2374) & _GEN_2342;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_14 <= ~(_GEN_2248 | _GEN_2375) & _GEN_2343;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_15 <= ~(_GEN_2249 | _GEN_2376) & _GEN_2344;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_16 <= ~(_GEN_2250 | _GEN_2377) & _GEN_2345;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_17 <= ~(_GEN_2251 | _GEN_2378) & _GEN_2346;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_18 <= ~(_GEN_2252 | _GEN_2379) & _GEN_2347;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_19 <= ~(_GEN_2253 | _GEN_2380) & _GEN_2348;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_20 <= ~(_GEN_2254 | _GEN_2381) & _GEN_2349;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_21 <= ~(_GEN_2255 | _GEN_2382) & _GEN_2350;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_22 <= ~(_GEN_2256 | _GEN_2383) & _GEN_2351;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_23 <= ~(_GEN_2257 | _GEN_2384) & _GEN_2352;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_24 <= ~(_GEN_2258 | _GEN_2385) & _GEN_2353;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_25 <= ~(_GEN_2259 | _GEN_2386) & _GEN_2354;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_26 <= ~(_GEN_2260 | _GEN_2387) & _GEN_2355;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_27 <= ~(_GEN_2261 | _GEN_2388) & _GEN_2356;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_28 <= ~(_GEN_2262 | _GEN_2389) & _GEN_2357;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_29 <= ~(_GEN_2263 | _GEN_2390) & _GEN_2358;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_30 <= ~(_GEN_2264 | _GEN_2391) & _GEN_2359;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
        rob_val_2_31 <= ~((&rob_head) | _GEN_2392) & _GEN_2360;	// rob.scala:224:29, :307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20, :476:25
      end
      else begin	// rob.scala:547:70
        rob_val_2_0 <= ~_GEN_2361 & _GEN_2329;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_1 <= ~_GEN_2362 & _GEN_2330;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_2 <= ~_GEN_2363 & _GEN_2331;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_3 <= ~_GEN_2364 & _GEN_2332;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_4 <= ~_GEN_2365 & _GEN_2333;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_5 <= ~_GEN_2366 & _GEN_2334;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_6 <= ~_GEN_2367 & _GEN_2335;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_7 <= ~_GEN_2368 & _GEN_2336;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_8 <= ~_GEN_2369 & _GEN_2337;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_9 <= ~_GEN_2370 & _GEN_2338;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_10 <= ~_GEN_2371 & _GEN_2339;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_11 <= ~_GEN_2372 & _GEN_2340;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_12 <= ~_GEN_2373 & _GEN_2341;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_13 <= ~_GEN_2374 & _GEN_2342;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_14 <= ~_GEN_2375 & _GEN_2343;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_15 <= ~_GEN_2376 & _GEN_2344;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_16 <= ~_GEN_2377 & _GEN_2345;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_17 <= ~_GEN_2378 & _GEN_2346;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_18 <= ~_GEN_2379 & _GEN_2347;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_19 <= ~_GEN_2380 & _GEN_2348;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_20 <= ~_GEN_2381 & _GEN_2349;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_21 <= ~_GEN_2382 & _GEN_2350;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_22 <= ~_GEN_2383 & _GEN_2351;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_23 <= ~_GEN_2384 & _GEN_2352;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_24 <= ~_GEN_2385 & _GEN_2353;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_25 <= ~_GEN_2386 & _GEN_2354;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_26 <= ~_GEN_2387 & _GEN_2355;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_27 <= ~_GEN_2388 & _GEN_2356;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_28 <= ~_GEN_2389 & _GEN_2357;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_29 <= ~_GEN_2390 & _GEN_2358;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_30 <= ~_GEN_2391 & _GEN_2359;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
        rob_val_2_31 <= ~_GEN_2392 & _GEN_2360;	// rob.scala:307:32, :323:29, :324:31, :433:20, :434:30, :455:7, :456:20
      end
      if (io_enq_valids_0 | io_enq_valids_1 | io_enq_valids_2)	// rob.scala:679:31
        r_partial_row <= io_enq_partial_stall;	// rob.scala:677:30
      pnr_maybe_at_tail <= ~rob_deq & (do_inc_row | pnr_maybe_at_tail);	// rob.scala:688:34, :714:36, :717:52, :736:{26,35,50}, :750:76, :754:13
    end
    r_xcpt_uop_br_mask <= next_xcpt_uop_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:259:29, :625:17, :631:76, :632:27, util.scala:85:{25,27}
    if (_GEN_2165) begin	// rob.scala:631:47
      if (io_lxcpt_valid) begin
        if (_GEN_2166) begin	// rob.scala:635:25
          r_xcpt_uop_rob_idx <= io_lxcpt_bits_uop_rob_idx;	// rob.scala:259:29
          r_xcpt_uop_exc_cause <= {59'h0, io_lxcpt_bits_cause};	// rob.scala:259:29, :556:50, :638:33
          r_xcpt_badvaddr <= io_lxcpt_bits_badvaddr;	// rob.scala:260:29
        end
      end
      else if (_GEN_2167) begin	// rob.scala:641:30
        automatic logic [3:0][6:0]  _GEN_2400 =
          {{io_enq_uops_0_rob_idx},
           {io_enq_uops_2_rob_idx},
           {io_enq_uops_1_rob_idx},
           {io_enq_uops_0_rob_idx}};	// rob.scala:646:23
        automatic logic [3:0][63:0] _GEN_2401 =
          {{io_enq_uops_0_exc_cause},
           {io_enq_uops_2_exc_cause},
           {io_enq_uops_1_exc_cause},
           {io_enq_uops_0_exc_cause}};	// rob.scala:646:23
        automatic logic [3:0][5:0]  _GEN_2402 =
          {{io_enq_uops_0_pc_lob},
           {io_enq_uops_2_pc_lob},
           {io_enq_uops_1_pc_lob},
           {io_enq_uops_0_pc_lob}};	// rob.scala:646:23
        r_xcpt_uop_rob_idx <= _GEN_2400[idx];	// rob.scala:259:29, :642:37, :646:23
        r_xcpt_uop_exc_cause <= _GEN_2401[idx];	// rob.scala:259:29, :642:37, :646:23
        r_xcpt_badvaddr <= {io_xcpt_fetch_pc[39:6], _GEN_2402[idx]};	// rob.scala:260:29, :642:37, :646:23, :647:76
      end
    end
    if (_GEN_8) begin	// rob.scala:361:31
      automatic logic _GEN_2403;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2404;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2405;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2406;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2407;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2408;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2409;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2410;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2411;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2412;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2413;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2414;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2415;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2416;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2417;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2418;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2419;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2420;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2421;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2422;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2423;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2424;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2425;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2426;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2427;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2428;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2429;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2430;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2431;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2432;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2433;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2434;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2403 = _GEN_856 | _GEN_794;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2404 = _GEN_857 | _GEN_796;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2405 = _GEN_858 | _GEN_798;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2406 = _GEN_859 | _GEN_800;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2407 = _GEN_860 | _GEN_802;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2408 = _GEN_861 | _GEN_804;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2409 = _GEN_862 | _GEN_806;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2410 = _GEN_863 | _GEN_808;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2411 = _GEN_864 | _GEN_810;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2412 = _GEN_865 | _GEN_812;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2413 = _GEN_866 | _GEN_814;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2414 = _GEN_867 | _GEN_816;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2415 = _GEN_868 | _GEN_818;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2416 = _GEN_869 | _GEN_820;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2417 = _GEN_870 | _GEN_822;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2418 = _GEN_871 | _GEN_824;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2419 = _GEN_872 | _GEN_826;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2420 = _GEN_873 | _GEN_828;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2421 = _GEN_874 | _GEN_830;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2422 = _GEN_875 | _GEN_832;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2423 = _GEN_876 | _GEN_834;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2424 = _GEN_877 | _GEN_836;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2425 = _GEN_878 | _GEN_838;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2426 = _GEN_879 | _GEN_840;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2427 = _GEN_880 | _GEN_842;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2428 = _GEN_881 | _GEN_844;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2429 = _GEN_882 | _GEN_846;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2430 = _GEN_883 | _GEN_848;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2431 = _GEN_884 | _GEN_850;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2432 = _GEN_885 | _GEN_852;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2433 = _GEN_886 | _GEN_854;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2434 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_855;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
      rob_bsy_0 <= ~_GEN_2403 & _GEN_668;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1 <= ~_GEN_2404 & _GEN_671;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2 <= ~_GEN_2405 & _GEN_674;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_3 <= ~_GEN_2406 & _GEN_677;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_4 <= ~_GEN_2407 & _GEN_680;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_5 <= ~_GEN_2408 & _GEN_683;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_6 <= ~_GEN_2409 & _GEN_686;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_7 <= ~_GEN_2410 & _GEN_689;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_8 <= ~_GEN_2411 & _GEN_692;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_9 <= ~_GEN_2412 & _GEN_695;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_10 <= ~_GEN_2413 & _GEN_698;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_11 <= ~_GEN_2414 & _GEN_701;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_12 <= ~_GEN_2415 & _GEN_704;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_13 <= ~_GEN_2416 & _GEN_707;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_14 <= ~_GEN_2417 & _GEN_710;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_15 <= ~_GEN_2418 & _GEN_713;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_16 <= ~_GEN_2419 & _GEN_716;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_17 <= ~_GEN_2420 & _GEN_719;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_18 <= ~_GEN_2421 & _GEN_722;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_19 <= ~_GEN_2422 & _GEN_725;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_20 <= ~_GEN_2423 & _GEN_728;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_21 <= ~_GEN_2424 & _GEN_731;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_22 <= ~_GEN_2425 & _GEN_734;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_23 <= ~_GEN_2426 & _GEN_737;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_24 <= ~_GEN_2427 & _GEN_740;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_25 <= ~_GEN_2428 & _GEN_743;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_26 <= ~_GEN_2429 & _GEN_746;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_27 <= ~_GEN_2430 & _GEN_749;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_28 <= ~_GEN_2431 & _GEN_752;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_29 <= ~_GEN_2432 & _GEN_755;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_30 <= ~_GEN_2433 & _GEN_758;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_31 <= ~_GEN_2434 & _GEN_760;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_unsafe_0 <= ~_GEN_2403 & _GEN_761;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1 <= ~_GEN_2404 & _GEN_762;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2 <= ~_GEN_2405 & _GEN_763;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_3 <= ~_GEN_2406 & _GEN_764;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_4 <= ~_GEN_2407 & _GEN_765;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_5 <= ~_GEN_2408 & _GEN_766;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_6 <= ~_GEN_2409 & _GEN_767;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_7 <= ~_GEN_2410 & _GEN_768;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_8 <= ~_GEN_2411 & _GEN_769;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_9 <= ~_GEN_2412 & _GEN_770;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_10 <= ~_GEN_2413 & _GEN_771;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_11 <= ~_GEN_2414 & _GEN_772;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_12 <= ~_GEN_2415 & _GEN_773;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_13 <= ~_GEN_2416 & _GEN_774;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_14 <= ~_GEN_2417 & _GEN_775;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_15 <= ~_GEN_2418 & _GEN_776;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_16 <= ~_GEN_2419 & _GEN_777;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_17 <= ~_GEN_2420 & _GEN_778;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_18 <= ~_GEN_2421 & _GEN_779;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_19 <= ~_GEN_2422 & _GEN_780;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_20 <= ~_GEN_2423 & _GEN_781;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_21 <= ~_GEN_2424 & _GEN_782;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_22 <= ~_GEN_2425 & _GEN_783;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_23 <= ~_GEN_2426 & _GEN_784;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_24 <= ~_GEN_2427 & _GEN_785;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_25 <= ~_GEN_2428 & _GEN_786;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_26 <= ~_GEN_2429 & _GEN_787;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_27 <= ~_GEN_2430 & _GEN_788;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_28 <= ~_GEN_2431 & _GEN_789;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_29 <= ~_GEN_2432 & _GEN_790;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_30 <= ~_GEN_2433 & _GEN_791;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_31 <= ~_GEN_2434 & _GEN_792;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
    end
    else begin	// rob.scala:361:31
      rob_bsy_0 <= ~_GEN_794 & _GEN_668;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1 <= ~_GEN_796 & _GEN_671;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2 <= ~_GEN_798 & _GEN_674;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_3 <= ~_GEN_800 & _GEN_677;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_4 <= ~_GEN_802 & _GEN_680;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_5 <= ~_GEN_804 & _GEN_683;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_6 <= ~_GEN_806 & _GEN_686;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_7 <= ~_GEN_808 & _GEN_689;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_8 <= ~_GEN_810 & _GEN_692;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_9 <= ~_GEN_812 & _GEN_695;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_10 <= ~_GEN_814 & _GEN_698;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_11 <= ~_GEN_816 & _GEN_701;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_12 <= ~_GEN_818 & _GEN_704;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_13 <= ~_GEN_820 & _GEN_707;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_14 <= ~_GEN_822 & _GEN_710;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_15 <= ~_GEN_824 & _GEN_713;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_16 <= ~_GEN_826 & _GEN_716;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_17 <= ~_GEN_828 & _GEN_719;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_18 <= ~_GEN_830 & _GEN_722;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_19 <= ~_GEN_832 & _GEN_725;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_20 <= ~_GEN_834 & _GEN_728;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_21 <= ~_GEN_836 & _GEN_731;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_22 <= ~_GEN_838 & _GEN_734;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_23 <= ~_GEN_840 & _GEN_737;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_24 <= ~_GEN_842 & _GEN_740;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_25 <= ~_GEN_844 & _GEN_743;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_26 <= ~_GEN_846 & _GEN_746;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_27 <= ~_GEN_848 & _GEN_749;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_28 <= ~_GEN_850 & _GEN_752;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_29 <= ~_GEN_852 & _GEN_755;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_30 <= ~_GEN_854 & _GEN_758;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_31 <= ~_GEN_855 & _GEN_760;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_unsafe_0 <= ~_GEN_794 & _GEN_761;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1 <= ~_GEN_796 & _GEN_762;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2 <= ~_GEN_798 & _GEN_763;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_3 <= ~_GEN_800 & _GEN_764;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_4 <= ~_GEN_802 & _GEN_765;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_5 <= ~_GEN_804 & _GEN_766;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_6 <= ~_GEN_806 & _GEN_767;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_7 <= ~_GEN_808 & _GEN_768;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_8 <= ~_GEN_810 & _GEN_769;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_9 <= ~_GEN_812 & _GEN_770;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_10 <= ~_GEN_814 & _GEN_771;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_11 <= ~_GEN_816 & _GEN_772;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_12 <= ~_GEN_818 & _GEN_773;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_13 <= ~_GEN_820 & _GEN_774;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_14 <= ~_GEN_822 & _GEN_775;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_15 <= ~_GEN_824 & _GEN_776;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_16 <= ~_GEN_826 & _GEN_777;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_17 <= ~_GEN_828 & _GEN_778;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_18 <= ~_GEN_830 & _GEN_779;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_19 <= ~_GEN_832 & _GEN_780;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_20 <= ~_GEN_834 & _GEN_781;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_21 <= ~_GEN_836 & _GEN_782;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_22 <= ~_GEN_838 & _GEN_783;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_23 <= ~_GEN_840 & _GEN_784;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_24 <= ~_GEN_842 & _GEN_785;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_25 <= ~_GEN_844 & _GEN_786;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_26 <= ~_GEN_846 & _GEN_787;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_27 <= ~_GEN_848 & _GEN_788;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_28 <= ~_GEN_850 & _GEN_789;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_29 <= ~_GEN_852 & _GEN_790;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_30 <= ~_GEN_854 & _GEN_791;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_31 <= ~_GEN_855 & _GEN_792;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
    end
    if (_GEN_97) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_0_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_0_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_0_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_0_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_0_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_0_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_0_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_0_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_0_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_0_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_0_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_0_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_0_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_0_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_0_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_0_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_981) | ~rob_val_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_97)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_0_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_0_br_mask <= rob_uop_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_99) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_1_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_1_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_1_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_1_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_1_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_1_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_1_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_1_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_1_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_1_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_1_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_1_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_1_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_982) | ~rob_val_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_99)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_br_mask <= rob_uop_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_101) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_2_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_2_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_2_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_2_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_2_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_2_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_2_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_2_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_2_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_2_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_2_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_2_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_2_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_983) | ~rob_val_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_101)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_br_mask <= rob_uop_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_103) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_3_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_3_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_3_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_3_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_3_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_3_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_3_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_3_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_3_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_3_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_3_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_3_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_3_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_3_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_3_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_3_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_984) | ~rob_val_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_103)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_3_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_3_br_mask <= rob_uop_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_105) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_4_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_4_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_4_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_4_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_4_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_4_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_4_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_4_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_4_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_4_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_4_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_4_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_4_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_4_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_4_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_4_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_985) | ~rob_val_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_105)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_4_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_4_br_mask <= rob_uop_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_107) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_5_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_5_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_5_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_5_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_5_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_5_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_5_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_5_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_5_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_5_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_5_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_5_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_5_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_5_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_5_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_5_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_986) | ~rob_val_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_107)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_5_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_5_br_mask <= rob_uop_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_109) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_6_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_6_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_6_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_6_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_6_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_6_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_6_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_6_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_6_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_6_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_6_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_6_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_6_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_6_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_6_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_6_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_987) | ~rob_val_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_109)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_6_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_6_br_mask <= rob_uop_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_111) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_7_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_7_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_7_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_7_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_7_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_7_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_7_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_7_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_7_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_7_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_7_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_7_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_7_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_7_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_7_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_7_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_988) | ~rob_val_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_111)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_7_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_7_br_mask <= rob_uop_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_113) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_8_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_8_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_8_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_8_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_8_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_8_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_8_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_8_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_8_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_8_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_8_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_8_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_8_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_8_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_8_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_8_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_989) | ~rob_val_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_113)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_8_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_8_br_mask <= rob_uop_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_115) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_9_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_9_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_9_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_9_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_9_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_9_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_9_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_9_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_9_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_9_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_9_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_9_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_9_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_9_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_9_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_9_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_990) | ~rob_val_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_115)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_9_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_9_br_mask <= rob_uop_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_117) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_10_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_10_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_10_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_10_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_10_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_10_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_10_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_10_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_10_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_10_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_10_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_10_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_10_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_10_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_10_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_10_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_991) | ~rob_val_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_117)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_10_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_10_br_mask <= rob_uop_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_119) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_11_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_11_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_11_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_11_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_11_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_11_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_11_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_11_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_11_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_11_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_11_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_11_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_11_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_11_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_11_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_11_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_992) | ~rob_val_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_119)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_11_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_11_br_mask <= rob_uop_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_121) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_12_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_12_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_12_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_12_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_12_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_12_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_12_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_12_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_12_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_12_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_12_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_12_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_12_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_12_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_12_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_12_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_993) | ~rob_val_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_121)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_12_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_12_br_mask <= rob_uop_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_123) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_13_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_13_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_13_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_13_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_13_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_13_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_13_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_13_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_13_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_13_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_13_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_13_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_13_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_13_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_13_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_13_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_994) | ~rob_val_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_123)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_13_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_13_br_mask <= rob_uop_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_125) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_14_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_14_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_14_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_14_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_14_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_14_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_14_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_14_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_14_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_14_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_14_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_14_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_14_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_14_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_14_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_14_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_995) | ~rob_val_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_125)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_14_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_14_br_mask <= rob_uop_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_127) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_15_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_15_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_15_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_15_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_15_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_15_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_15_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_15_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_15_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_15_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_15_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_15_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_15_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_15_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_15_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_15_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_996) | ~rob_val_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_127)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_15_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_15_br_mask <= rob_uop_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_129) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_16_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_16_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_16_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_16_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_16_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_16_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_16_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_16_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_16_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_16_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_16_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_16_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_16_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_16_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_16_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_16_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_997) | ~rob_val_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_129)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_16_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_16_br_mask <= rob_uop_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_131) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_17_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_17_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_17_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_17_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_17_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_17_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_17_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_17_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_17_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_17_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_17_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_17_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_17_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_17_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_17_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_17_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_998) | ~rob_val_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_131)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_17_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_17_br_mask <= rob_uop_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_133) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_18_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_18_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_18_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_18_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_18_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_18_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_18_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_18_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_18_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_18_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_18_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_18_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_18_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_18_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_18_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_18_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_999) | ~rob_val_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_133)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_18_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_18_br_mask <= rob_uop_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_135) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_19_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_19_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_19_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_19_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_19_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_19_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_19_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_19_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_19_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_19_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_19_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_19_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_19_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_19_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_19_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_19_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1000) | ~rob_val_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_135)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_19_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_19_br_mask <= rob_uop_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_137) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_20_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_20_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_20_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_20_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_20_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_20_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_20_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_20_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_20_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_20_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_20_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_20_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_20_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_20_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_20_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_20_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1001) | ~rob_val_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_137)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_20_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_20_br_mask <= rob_uop_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_139) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_21_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_21_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_21_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_21_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_21_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_21_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_21_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_21_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_21_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_21_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_21_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_21_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_21_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_21_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_21_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_21_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1002) | ~rob_val_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_139)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_21_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_21_br_mask <= rob_uop_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_141) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_22_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_22_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_22_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_22_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_22_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_22_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_22_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_22_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_22_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_22_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_22_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_22_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_22_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_22_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_22_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_22_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1003) | ~rob_val_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_141)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_22_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_22_br_mask <= rob_uop_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_143) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_23_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_23_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_23_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_23_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_23_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_23_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_23_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_23_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_23_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_23_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_23_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_23_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_23_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_23_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_23_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_23_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1004) | ~rob_val_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_143)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_23_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_23_br_mask <= rob_uop_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_145) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_24_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_24_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_24_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_24_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_24_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_24_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_24_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_24_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_24_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_24_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_24_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_24_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_24_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_24_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_24_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_24_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1005) | ~rob_val_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_145)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_24_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_24_br_mask <= rob_uop_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_147) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_25_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_25_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_25_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_25_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_25_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_25_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_25_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_25_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_25_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_25_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_25_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_25_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_25_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_25_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_25_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_25_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1006) | ~rob_val_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_147)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_25_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_25_br_mask <= rob_uop_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_149) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_26_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_26_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_26_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_26_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_26_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_26_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_26_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_26_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_26_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_26_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_26_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_26_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_26_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_26_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_26_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_26_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1007) | ~rob_val_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_149)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_26_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_26_br_mask <= rob_uop_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_151) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_27_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_27_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_27_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_27_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_27_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_27_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_27_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_27_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_27_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_27_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_27_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_27_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_27_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_27_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_27_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_27_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1008) | ~rob_val_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_151)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_27_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_27_br_mask <= rob_uop_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_153) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_28_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_28_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_28_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_28_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_28_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_28_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_28_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_28_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_28_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_28_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_28_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_28_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_28_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_28_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_28_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_28_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1009) | ~rob_val_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_153)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_28_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_28_br_mask <= rob_uop_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_155) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_29_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_29_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_29_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_29_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_29_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_29_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_29_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_29_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_29_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_29_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_29_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_29_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_29_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_29_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_29_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_29_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1010) | ~rob_val_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_155)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_29_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_29_br_mask <= rob_uop_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_157) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_30_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_30_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_30_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_30_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_30_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_30_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_30_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_30_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_30_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_30_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_30_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_30_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_30_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_30_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_30_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_30_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1011) | ~rob_val_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_157)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_30_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_30_br_mask <= rob_uop_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_158) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_31_uopc <= io_enq_uops_0_uopc;	// rob.scala:310:28
      rob_uop_31_is_rvc <= io_enq_uops_0_is_rvc;	// rob.scala:310:28
      rob_uop_31_ftq_idx <= io_enq_uops_0_ftq_idx;	// rob.scala:310:28
      rob_uop_31_edge_inst <= io_enq_uops_0_edge_inst;	// rob.scala:310:28
      rob_uop_31_pc_lob <= io_enq_uops_0_pc_lob;	// rob.scala:310:28
      rob_uop_31_pdst <= io_enq_uops_0_pdst;	// rob.scala:310:28
      rob_uop_31_stale_pdst <= io_enq_uops_0_stale_pdst;	// rob.scala:310:28
      rob_uop_31_is_fencei <= io_enq_uops_0_is_fencei;	// rob.scala:310:28
      rob_uop_31_uses_ldq <= io_enq_uops_0_uses_ldq;	// rob.scala:310:28
      rob_uop_31_uses_stq <= io_enq_uops_0_uses_stq;	// rob.scala:310:28
      rob_uop_31_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_31_flush_on_commit <= io_enq_uops_0_flush_on_commit;	// rob.scala:310:28
      rob_uop_31_ldst <= io_enq_uops_0_ldst;	// rob.scala:310:28
      rob_uop_31_ldst_val <= io_enq_uops_0_ldst_val;	// rob.scala:310:28
      rob_uop_31_dst_rtype <= io_enq_uops_0_dst_rtype;	// rob.scala:310:28
      rob_uop_31_fp_val <= io_enq_uops_0_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1012) | ~rob_val_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_158)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_31_br_mask <= io_enq_uops_0_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_31_br_mask <= rob_uop_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_0 <=
      ~_GEN_919
      & (_GEN_9 & _GEN_887 | (_GEN_97 ? io_enq_uops_0_exception : rob_exception_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1 <=
      ~_GEN_921
      & (_GEN_9 & _GEN_888 | (_GEN_99 ? io_enq_uops_0_exception : rob_exception_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2 <=
      ~_GEN_923
      & (_GEN_9 & _GEN_889 | (_GEN_101 ? io_enq_uops_0_exception : rob_exception_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_3 <=
      ~_GEN_925
      & (_GEN_9 & _GEN_890 | (_GEN_103 ? io_enq_uops_0_exception : rob_exception_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_4 <=
      ~_GEN_927
      & (_GEN_9 & _GEN_891 | (_GEN_105 ? io_enq_uops_0_exception : rob_exception_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_5 <=
      ~_GEN_929
      & (_GEN_9 & _GEN_892 | (_GEN_107 ? io_enq_uops_0_exception : rob_exception_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_6 <=
      ~_GEN_931
      & (_GEN_9 & _GEN_893 | (_GEN_109 ? io_enq_uops_0_exception : rob_exception_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_7 <=
      ~_GEN_933
      & (_GEN_9 & _GEN_894 | (_GEN_111 ? io_enq_uops_0_exception : rob_exception_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_8 <=
      ~_GEN_935
      & (_GEN_9 & _GEN_895 | (_GEN_113 ? io_enq_uops_0_exception : rob_exception_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_9 <=
      ~_GEN_937
      & (_GEN_9 & _GEN_896 | (_GEN_115 ? io_enq_uops_0_exception : rob_exception_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_10 <=
      ~_GEN_939
      & (_GEN_9 & _GEN_897 | (_GEN_117 ? io_enq_uops_0_exception : rob_exception_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_11 <=
      ~_GEN_941
      & (_GEN_9 & _GEN_898 | (_GEN_119 ? io_enq_uops_0_exception : rob_exception_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_12 <=
      ~_GEN_943
      & (_GEN_9 & _GEN_899 | (_GEN_121 ? io_enq_uops_0_exception : rob_exception_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_13 <=
      ~_GEN_945
      & (_GEN_9 & _GEN_900 | (_GEN_123 ? io_enq_uops_0_exception : rob_exception_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_14 <=
      ~_GEN_947
      & (_GEN_9 & _GEN_901 | (_GEN_125 ? io_enq_uops_0_exception : rob_exception_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_15 <=
      ~_GEN_949
      & (_GEN_9 & _GEN_902 | (_GEN_127 ? io_enq_uops_0_exception : rob_exception_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_16 <=
      ~_GEN_951
      & (_GEN_9 & _GEN_903 | (_GEN_129 ? io_enq_uops_0_exception : rob_exception_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_17 <=
      ~_GEN_953
      & (_GEN_9 & _GEN_904 | (_GEN_131 ? io_enq_uops_0_exception : rob_exception_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_18 <=
      ~_GEN_955
      & (_GEN_9 & _GEN_905 | (_GEN_133 ? io_enq_uops_0_exception : rob_exception_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_19 <=
      ~_GEN_957
      & (_GEN_9 & _GEN_906 | (_GEN_135 ? io_enq_uops_0_exception : rob_exception_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_20 <=
      ~_GEN_959
      & (_GEN_9 & _GEN_907 | (_GEN_137 ? io_enq_uops_0_exception : rob_exception_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_21 <=
      ~_GEN_961
      & (_GEN_9 & _GEN_908 | (_GEN_139 ? io_enq_uops_0_exception : rob_exception_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_22 <=
      ~_GEN_963
      & (_GEN_9 & _GEN_909 | (_GEN_141 ? io_enq_uops_0_exception : rob_exception_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_23 <=
      ~_GEN_965
      & (_GEN_9 & _GEN_910 | (_GEN_143 ? io_enq_uops_0_exception : rob_exception_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_24 <=
      ~_GEN_967
      & (_GEN_9 & _GEN_911 | (_GEN_145 ? io_enq_uops_0_exception : rob_exception_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_25 <=
      ~_GEN_969
      & (_GEN_9 & _GEN_912 | (_GEN_147 ? io_enq_uops_0_exception : rob_exception_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_26 <=
      ~_GEN_971
      & (_GEN_9 & _GEN_913 | (_GEN_149 ? io_enq_uops_0_exception : rob_exception_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_27 <=
      ~_GEN_973
      & (_GEN_9 & _GEN_914 | (_GEN_151 ? io_enq_uops_0_exception : rob_exception_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_28 <=
      ~_GEN_975
      & (_GEN_9 & _GEN_915 | (_GEN_153 ? io_enq_uops_0_exception : rob_exception_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_29 <=
      ~_GEN_977
      & (_GEN_9 & _GEN_916 | (_GEN_155 ? io_enq_uops_0_exception : rob_exception_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_30 <=
      ~_GEN_979
      & (_GEN_9 & _GEN_917 | (_GEN_157 ? io_enq_uops_0_exception : rob_exception_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_31 <=
      ~_GEN_980
      & (_GEN_9 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_158 ? io_enq_uops_0_exception : rob_exception_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_0 <=
      ~(_GEN_5 & _GEN_666)
      & (_GEN_604
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_476 | _GEN_414 | _GEN_1 & _GEN_286)
             & (_GEN_224 ? io_wb_resps_0_bits_predicated : ~_GEN_97 & rob_predicated_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1 <=
      ~(_GEN_5 & _GEN_669)
      & (_GEN_606
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_479 | _GEN_416 | _GEN_1 & _GEN_289)
             & (_GEN_226 ? io_wb_resps_0_bits_predicated : ~_GEN_99 & rob_predicated_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2 <=
      ~(_GEN_5 & _GEN_672)
      & (_GEN_608
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_482 | _GEN_418 | _GEN_1 & _GEN_292)
             & (_GEN_228 ? io_wb_resps_0_bits_predicated : ~_GEN_101 & rob_predicated_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_3 <=
      ~(_GEN_5 & _GEN_675)
      & (_GEN_610
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_485 | _GEN_420 | _GEN_1 & _GEN_295)
             & (_GEN_230 ? io_wb_resps_0_bits_predicated : ~_GEN_103 & rob_predicated_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_4 <=
      ~(_GEN_5 & _GEN_678)
      & (_GEN_612
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_488 | _GEN_422 | _GEN_1 & _GEN_298)
             & (_GEN_232 ? io_wb_resps_0_bits_predicated : ~_GEN_105 & rob_predicated_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_5 <=
      ~(_GEN_5 & _GEN_681)
      & (_GEN_614
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_491 | _GEN_424 | _GEN_1 & _GEN_301)
             & (_GEN_234 ? io_wb_resps_0_bits_predicated : ~_GEN_107 & rob_predicated_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_6 <=
      ~(_GEN_5 & _GEN_684)
      & (_GEN_616
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_494 | _GEN_426 | _GEN_1 & _GEN_304)
             & (_GEN_236 ? io_wb_resps_0_bits_predicated : ~_GEN_109 & rob_predicated_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_7 <=
      ~(_GEN_5 & _GEN_687)
      & (_GEN_618
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_497 | _GEN_428 | _GEN_1 & _GEN_307)
             & (_GEN_238 ? io_wb_resps_0_bits_predicated : ~_GEN_111 & rob_predicated_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_8 <=
      ~(_GEN_5 & _GEN_690)
      & (_GEN_620
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_500 | _GEN_430 | _GEN_1 & _GEN_310)
             & (_GEN_240 ? io_wb_resps_0_bits_predicated : ~_GEN_113 & rob_predicated_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_9 <=
      ~(_GEN_5 & _GEN_693)
      & (_GEN_622
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_503 | _GEN_432 | _GEN_1 & _GEN_313)
             & (_GEN_242 ? io_wb_resps_0_bits_predicated : ~_GEN_115 & rob_predicated_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_10 <=
      ~(_GEN_5 & _GEN_696)
      & (_GEN_624
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_506 | _GEN_434 | _GEN_1 & _GEN_316)
             & (_GEN_244
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_117 & rob_predicated_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_11 <=
      ~(_GEN_5 & _GEN_699)
      & (_GEN_626
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_509 | _GEN_436 | _GEN_1 & _GEN_319)
             & (_GEN_246
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_119 & rob_predicated_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_12 <=
      ~(_GEN_5 & _GEN_702)
      & (_GEN_628
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_512 | _GEN_438 | _GEN_1 & _GEN_322)
             & (_GEN_248
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_121 & rob_predicated_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_13 <=
      ~(_GEN_5 & _GEN_705)
      & (_GEN_630
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_515 | _GEN_440 | _GEN_1 & _GEN_325)
             & (_GEN_250
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_123 & rob_predicated_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_14 <=
      ~(_GEN_5 & _GEN_708)
      & (_GEN_632
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_518 | _GEN_442 | _GEN_1 & _GEN_328)
             & (_GEN_252
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_125 & rob_predicated_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_15 <=
      ~(_GEN_5 & _GEN_711)
      & (_GEN_634
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_521 | _GEN_444 | _GEN_1 & _GEN_331)
             & (_GEN_254
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_127 & rob_predicated_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_16 <=
      ~(_GEN_5 & _GEN_714)
      & (_GEN_636
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_524 | _GEN_446 | _GEN_1 & _GEN_334)
             & (_GEN_256
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_129 & rob_predicated_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_17 <=
      ~(_GEN_5 & _GEN_717)
      & (_GEN_638
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_527 | _GEN_448 | _GEN_1 & _GEN_337)
             & (_GEN_258
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_131 & rob_predicated_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_18 <=
      ~(_GEN_5 & _GEN_720)
      & (_GEN_640
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_530 | _GEN_450 | _GEN_1 & _GEN_340)
             & (_GEN_260
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_133 & rob_predicated_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_19 <=
      ~(_GEN_5 & _GEN_723)
      & (_GEN_642
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_533 | _GEN_452 | _GEN_1 & _GEN_343)
             & (_GEN_262
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_135 & rob_predicated_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_20 <=
      ~(_GEN_5 & _GEN_726)
      & (_GEN_644
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_536 | _GEN_454 | _GEN_1 & _GEN_346)
             & (_GEN_264
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_137 & rob_predicated_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_21 <=
      ~(_GEN_5 & _GEN_729)
      & (_GEN_646
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_539 | _GEN_456 | _GEN_1 & _GEN_349)
             & (_GEN_266
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_139 & rob_predicated_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_22 <=
      ~(_GEN_5 & _GEN_732)
      & (_GEN_648
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_542 | _GEN_458 | _GEN_1 & _GEN_352)
             & (_GEN_268
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_141 & rob_predicated_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_23 <=
      ~(_GEN_5 & _GEN_735)
      & (_GEN_650
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_545 | _GEN_460 | _GEN_1 & _GEN_355)
             & (_GEN_270
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_143 & rob_predicated_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_24 <=
      ~(_GEN_5 & _GEN_738)
      & (_GEN_652
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_548 | _GEN_462 | _GEN_1 & _GEN_358)
             & (_GEN_272
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_145 & rob_predicated_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_25 <=
      ~(_GEN_5 & _GEN_741)
      & (_GEN_654
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_551 | _GEN_464 | _GEN_1 & _GEN_361)
             & (_GEN_274
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_147 & rob_predicated_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_26 <=
      ~(_GEN_5 & _GEN_744)
      & (_GEN_656
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_554 | _GEN_466 | _GEN_1 & _GEN_364)
             & (_GEN_276
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_149 & rob_predicated_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_27 <=
      ~(_GEN_5 & _GEN_747)
      & (_GEN_658
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_557 | _GEN_468 | _GEN_1 & _GEN_367)
             & (_GEN_278
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_151 & rob_predicated_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_28 <=
      ~(_GEN_5 & _GEN_750)
      & (_GEN_660
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_560 | _GEN_470 | _GEN_1 & _GEN_370)
             & (_GEN_280
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_153 & rob_predicated_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_29 <=
      ~(_GEN_5 & _GEN_753)
      & (_GEN_662
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_563 | _GEN_472 | _GEN_1 & _GEN_373)
             & (_GEN_282
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_155 & rob_predicated_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_30 <=
      ~(_GEN_5 & _GEN_756)
      & (_GEN_664
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & _GEN_566 | _GEN_474 | _GEN_1 & _GEN_376)
             & (_GEN_284
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_157 & rob_predicated_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_31 <=
      ~(_GEN_5 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])))
      & (_GEN_665
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_3 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_475 | _GEN_1
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_285
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_158 & rob_predicated_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    if (_GEN_38) begin	// rob.scala:361:31
      automatic logic _GEN_2435;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2436;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2437;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2438;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2439;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2440;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2441;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2442;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2443;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2444;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2445;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2446;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2447;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2448;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2449;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2450;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2451;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2452;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2453;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2454;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2455;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2456;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2457;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2458;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2459;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2460;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2461;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2462;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2463;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2464;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2465;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2466;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2435 = _GEN_856 | _GEN_1493;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2436 = _GEN_857 | _GEN_1494;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2437 = _GEN_858 | _GEN_1495;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2438 = _GEN_859 | _GEN_1496;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2439 = _GEN_860 | _GEN_1497;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2440 = _GEN_861 | _GEN_1498;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2441 = _GEN_862 | _GEN_1499;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2442 = _GEN_863 | _GEN_1500;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2443 = _GEN_864 | _GEN_1501;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2444 = _GEN_865 | _GEN_1502;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2445 = _GEN_866 | _GEN_1503;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2446 = _GEN_867 | _GEN_1504;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2447 = _GEN_868 | _GEN_1505;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2448 = _GEN_869 | _GEN_1506;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2449 = _GEN_870 | _GEN_1507;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2450 = _GEN_871 | _GEN_1508;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2451 = _GEN_872 | _GEN_1509;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2452 = _GEN_873 | _GEN_1510;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2453 = _GEN_874 | _GEN_1511;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2454 = _GEN_875 | _GEN_1512;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2455 = _GEN_876 | _GEN_1513;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2456 = _GEN_877 | _GEN_1514;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2457 = _GEN_878 | _GEN_1515;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2458 = _GEN_879 | _GEN_1516;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2459 = _GEN_880 | _GEN_1517;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2460 = _GEN_881 | _GEN_1518;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2461 = _GEN_882 | _GEN_1519;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2462 = _GEN_883 | _GEN_1520;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2463 = _GEN_884 | _GEN_1521;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2464 = _GEN_885 | _GEN_1522;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2465 = _GEN_886 | _GEN_1523;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2466 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_1524;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
      rob_bsy_1_0 <= ~_GEN_2435 & _GEN_1398;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_1 <= ~_GEN_2436 & _GEN_1400;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_2 <= ~_GEN_2437 & _GEN_1402;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_3 <= ~_GEN_2438 & _GEN_1404;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_4 <= ~_GEN_2439 & _GEN_1406;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_5 <= ~_GEN_2440 & _GEN_1408;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_6 <= ~_GEN_2441 & _GEN_1410;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_7 <= ~_GEN_2442 & _GEN_1412;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_8 <= ~_GEN_2443 & _GEN_1414;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_9 <= ~_GEN_2444 & _GEN_1416;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_10 <= ~_GEN_2445 & _GEN_1418;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_11 <= ~_GEN_2446 & _GEN_1420;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_12 <= ~_GEN_2447 & _GEN_1422;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_13 <= ~_GEN_2448 & _GEN_1424;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_14 <= ~_GEN_2449 & _GEN_1426;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_15 <= ~_GEN_2450 & _GEN_1428;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_16 <= ~_GEN_2451 & _GEN_1430;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_17 <= ~_GEN_2452 & _GEN_1432;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_18 <= ~_GEN_2453 & _GEN_1434;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_19 <= ~_GEN_2454 & _GEN_1436;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_20 <= ~_GEN_2455 & _GEN_1438;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_21 <= ~_GEN_2456 & _GEN_1440;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_22 <= ~_GEN_2457 & _GEN_1442;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_23 <= ~_GEN_2458 & _GEN_1444;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_24 <= ~_GEN_2459 & _GEN_1446;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_25 <= ~_GEN_2460 & _GEN_1448;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_26 <= ~_GEN_2461 & _GEN_1450;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_27 <= ~_GEN_2462 & _GEN_1452;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_28 <= ~_GEN_2463 & _GEN_1454;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_29 <= ~_GEN_2464 & _GEN_1456;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_30 <= ~_GEN_2465 & _GEN_1458;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_31 <= ~_GEN_2466 & _GEN_1460;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_unsafe_1_0 <= ~_GEN_2435 & _GEN_1461;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_1 <= ~_GEN_2436 & _GEN_1462;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_2 <= ~_GEN_2437 & _GEN_1463;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_3 <= ~_GEN_2438 & _GEN_1464;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_4 <= ~_GEN_2439 & _GEN_1465;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_5 <= ~_GEN_2440 & _GEN_1466;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_6 <= ~_GEN_2441 & _GEN_1467;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_7 <= ~_GEN_2442 & _GEN_1468;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_8 <= ~_GEN_2443 & _GEN_1469;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_9 <= ~_GEN_2444 & _GEN_1470;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_10 <= ~_GEN_2445 & _GEN_1471;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_11 <= ~_GEN_2446 & _GEN_1472;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_12 <= ~_GEN_2447 & _GEN_1473;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_13 <= ~_GEN_2448 & _GEN_1474;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_14 <= ~_GEN_2449 & _GEN_1475;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_15 <= ~_GEN_2450 & _GEN_1476;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_16 <= ~_GEN_2451 & _GEN_1477;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_17 <= ~_GEN_2452 & _GEN_1478;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_18 <= ~_GEN_2453 & _GEN_1479;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_19 <= ~_GEN_2454 & _GEN_1480;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_20 <= ~_GEN_2455 & _GEN_1481;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_21 <= ~_GEN_2456 & _GEN_1482;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_22 <= ~_GEN_2457 & _GEN_1483;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_23 <= ~_GEN_2458 & _GEN_1484;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_24 <= ~_GEN_2459 & _GEN_1485;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_25 <= ~_GEN_2460 & _GEN_1486;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_26 <= ~_GEN_2461 & _GEN_1487;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_27 <= ~_GEN_2462 & _GEN_1488;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_28 <= ~_GEN_2463 & _GEN_1489;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_29 <= ~_GEN_2464 & _GEN_1490;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_30 <= ~_GEN_2465 & _GEN_1491;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_31 <= ~_GEN_2466 & _GEN_1492;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
    end
    else begin	// rob.scala:361:31
      rob_bsy_1_0 <= ~_GEN_1493 & _GEN_1398;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_1 <= ~_GEN_1494 & _GEN_1400;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_2 <= ~_GEN_1495 & _GEN_1402;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_3 <= ~_GEN_1496 & _GEN_1404;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_4 <= ~_GEN_1497 & _GEN_1406;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_5 <= ~_GEN_1498 & _GEN_1408;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_6 <= ~_GEN_1499 & _GEN_1410;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_7 <= ~_GEN_1500 & _GEN_1412;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_8 <= ~_GEN_1501 & _GEN_1414;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_9 <= ~_GEN_1502 & _GEN_1416;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_10 <= ~_GEN_1503 & _GEN_1418;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_11 <= ~_GEN_1504 & _GEN_1420;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_12 <= ~_GEN_1505 & _GEN_1422;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_13 <= ~_GEN_1506 & _GEN_1424;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_14 <= ~_GEN_1507 & _GEN_1426;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_15 <= ~_GEN_1508 & _GEN_1428;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_16 <= ~_GEN_1509 & _GEN_1430;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_17 <= ~_GEN_1510 & _GEN_1432;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_18 <= ~_GEN_1511 & _GEN_1434;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_19 <= ~_GEN_1512 & _GEN_1436;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_20 <= ~_GEN_1513 & _GEN_1438;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_21 <= ~_GEN_1514 & _GEN_1440;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_22 <= ~_GEN_1515 & _GEN_1442;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_23 <= ~_GEN_1516 & _GEN_1444;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_24 <= ~_GEN_1517 & _GEN_1446;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_25 <= ~_GEN_1518 & _GEN_1448;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_26 <= ~_GEN_1519 & _GEN_1450;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_27 <= ~_GEN_1520 & _GEN_1452;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_28 <= ~_GEN_1521 & _GEN_1454;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_29 <= ~_GEN_1522 & _GEN_1456;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_30 <= ~_GEN_1523 & _GEN_1458;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_1_31 <= ~_GEN_1524 & _GEN_1460;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_unsafe_1_0 <= ~_GEN_1493 & _GEN_1461;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_1 <= ~_GEN_1494 & _GEN_1462;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_2 <= ~_GEN_1495 & _GEN_1463;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_3 <= ~_GEN_1496 & _GEN_1464;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_4 <= ~_GEN_1497 & _GEN_1465;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_5 <= ~_GEN_1498 & _GEN_1466;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_6 <= ~_GEN_1499 & _GEN_1467;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_7 <= ~_GEN_1500 & _GEN_1468;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_8 <= ~_GEN_1501 & _GEN_1469;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_9 <= ~_GEN_1502 & _GEN_1470;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_10 <= ~_GEN_1503 & _GEN_1471;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_11 <= ~_GEN_1504 & _GEN_1472;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_12 <= ~_GEN_1505 & _GEN_1473;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_13 <= ~_GEN_1506 & _GEN_1474;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_14 <= ~_GEN_1507 & _GEN_1475;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_15 <= ~_GEN_1508 & _GEN_1476;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_16 <= ~_GEN_1509 & _GEN_1477;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_17 <= ~_GEN_1510 & _GEN_1478;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_18 <= ~_GEN_1511 & _GEN_1479;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_19 <= ~_GEN_1512 & _GEN_1480;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_20 <= ~_GEN_1513 & _GEN_1481;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_21 <= ~_GEN_1514 & _GEN_1482;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_22 <= ~_GEN_1515 & _GEN_1483;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_23 <= ~_GEN_1516 & _GEN_1484;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_24 <= ~_GEN_1517 & _GEN_1485;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_25 <= ~_GEN_1518 & _GEN_1486;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_26 <= ~_GEN_1519 & _GEN_1487;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_27 <= ~_GEN_1520 & _GEN_1488;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_28 <= ~_GEN_1521 & _GEN_1489;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_29 <= ~_GEN_1522 & _GEN_1490;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_30 <= ~_GEN_1523 & _GEN_1491;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_1_31 <= ~_GEN_1524 & _GEN_1492;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
    end
    if (_GEN_1013) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_0_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_0_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_0_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_0_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_0_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_0_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_0_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_0_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_0_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_0_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_0_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_0_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_0_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_0_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_0_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_0_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1557) | ~rob_val_1_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1013)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_0_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_0_br_mask <= rob_uop_1_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1014) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_1_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_1_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_1_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_1_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_1_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_1_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_1_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_1_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_1_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_1_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_1_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_1_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_1_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_1_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_1_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_1_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1558) | ~rob_val_1_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1014)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_1_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_1_br_mask <= rob_uop_1_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1015) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_2_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_2_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_2_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_2_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_2_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_2_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_2_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_2_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_2_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_2_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_2_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_2_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_2_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_2_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_2_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_2_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1559) | ~rob_val_1_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1015)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_2_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_2_br_mask <= rob_uop_1_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1016) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_3_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_3_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_3_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_3_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_3_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_3_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_3_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_3_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_3_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_3_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_3_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_3_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_3_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_3_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_3_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_3_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1560) | ~rob_val_1_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1016)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_3_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_3_br_mask <= rob_uop_1_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1017) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_4_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_4_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_4_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_4_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_4_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_4_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_4_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_4_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_4_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_4_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_4_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_4_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_4_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_4_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_4_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_4_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1561) | ~rob_val_1_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1017)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_4_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_4_br_mask <= rob_uop_1_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1018) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_5_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_5_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_5_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_5_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_5_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_5_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_5_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_5_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_5_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_5_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_5_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_5_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_5_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_5_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_5_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_5_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1562) | ~rob_val_1_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1018)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_5_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_5_br_mask <= rob_uop_1_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1019) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_6_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_6_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_6_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_6_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_6_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_6_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_6_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_6_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_6_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_6_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_6_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_6_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_6_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_6_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_6_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_6_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1563) | ~rob_val_1_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1019)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_6_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_6_br_mask <= rob_uop_1_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1020) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_7_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_7_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_7_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_7_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_7_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_7_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_7_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_7_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_7_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_7_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_7_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_7_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_7_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_7_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_7_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_7_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1564) | ~rob_val_1_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1020)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_7_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_7_br_mask <= rob_uop_1_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1021) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_8_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_8_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_8_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_8_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_8_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_8_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_8_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_8_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_8_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_8_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_8_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_8_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_8_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_8_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_8_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_8_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1565) | ~rob_val_1_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1021)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_8_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_8_br_mask <= rob_uop_1_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1022) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_9_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_9_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_9_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_9_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_9_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_9_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_9_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_9_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_9_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_9_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_9_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_9_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_9_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_9_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_9_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_9_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1566) | ~rob_val_1_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1022)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_9_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_9_br_mask <= rob_uop_1_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1023) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_10_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_10_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_10_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_10_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_10_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_10_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_10_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_10_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_10_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_10_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_10_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_10_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_10_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_10_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_10_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_10_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1567) | ~rob_val_1_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1023)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_10_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_10_br_mask <= rob_uop_1_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1024) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_11_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_11_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_11_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_11_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_11_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_11_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_11_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_11_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_11_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_11_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_11_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_11_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_11_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_11_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_11_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_11_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1568) | ~rob_val_1_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1024)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_11_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_11_br_mask <= rob_uop_1_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1025) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_12_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_12_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_12_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_12_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_12_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_12_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_12_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_12_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_12_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_12_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_12_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_12_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_12_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_12_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_12_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_12_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1569) | ~rob_val_1_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1025)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_12_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_12_br_mask <= rob_uop_1_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1026) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_13_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_13_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_13_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_13_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_13_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_13_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_13_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_13_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_13_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_13_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_13_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_13_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_13_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_13_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_13_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_13_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1570) | ~rob_val_1_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1026)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_13_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_13_br_mask <= rob_uop_1_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1027) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_14_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_14_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_14_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_14_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_14_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_14_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_14_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_14_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_14_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_14_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_14_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_14_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_14_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_14_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_14_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_14_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1571) | ~rob_val_1_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1027)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_14_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_14_br_mask <= rob_uop_1_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1028) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_15_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_15_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_15_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_15_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_15_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_15_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_15_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_15_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_15_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_15_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_15_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_15_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_15_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_15_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_15_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_15_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1572) | ~rob_val_1_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1028)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_15_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_15_br_mask <= rob_uop_1_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1029) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_16_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_16_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_16_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_16_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_16_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_16_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_16_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_16_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_16_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_16_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_16_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_16_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_16_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_16_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_16_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_16_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1573) | ~rob_val_1_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1029)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_16_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_16_br_mask <= rob_uop_1_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1030) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_17_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_17_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_17_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_17_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_17_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_17_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_17_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_17_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_17_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_17_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_17_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_17_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_17_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_17_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_17_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_17_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1574) | ~rob_val_1_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1030)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_17_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_17_br_mask <= rob_uop_1_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1031) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_18_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_18_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_18_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_18_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_18_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_18_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_18_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_18_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_18_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_18_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_18_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_18_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_18_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_18_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_18_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_18_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1575) | ~rob_val_1_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1031)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_18_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_18_br_mask <= rob_uop_1_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1032) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_19_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_19_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_19_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_19_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_19_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_19_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_19_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_19_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_19_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_19_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_19_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_19_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_19_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_19_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_19_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_19_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1576) | ~rob_val_1_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1032)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_19_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_19_br_mask <= rob_uop_1_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1033) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_20_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_20_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_20_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_20_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_20_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_20_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_20_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_20_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_20_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_20_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_20_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_20_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_20_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_20_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_20_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_20_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1577) | ~rob_val_1_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1033)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_20_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_20_br_mask <= rob_uop_1_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1034) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_21_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_21_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_21_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_21_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_21_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_21_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_21_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_21_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_21_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_21_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_21_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_21_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_21_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_21_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_21_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_21_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1578) | ~rob_val_1_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1034)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_21_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_21_br_mask <= rob_uop_1_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1035) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_22_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_22_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_22_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_22_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_22_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_22_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_22_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_22_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_22_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_22_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_22_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_22_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_22_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_22_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_22_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_22_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1579) | ~rob_val_1_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1035)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_22_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_22_br_mask <= rob_uop_1_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1036) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_23_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_23_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_23_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_23_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_23_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_23_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_23_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_23_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_23_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_23_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_23_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_23_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_23_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_23_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_23_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_23_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1580) | ~rob_val_1_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1036)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_23_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_23_br_mask <= rob_uop_1_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1037) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_24_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_24_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_24_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_24_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_24_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_24_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_24_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_24_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_24_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_24_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_24_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_24_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_24_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_24_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_24_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_24_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1581) | ~rob_val_1_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1037)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_24_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_24_br_mask <= rob_uop_1_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1038) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_25_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_25_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_25_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_25_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_25_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_25_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_25_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_25_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_25_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_25_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_25_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_25_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_25_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_25_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_25_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_25_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1582) | ~rob_val_1_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1038)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_25_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_25_br_mask <= rob_uop_1_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1039) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_26_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_26_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_26_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_26_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_26_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_26_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_26_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_26_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_26_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_26_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_26_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_26_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_26_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_26_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_26_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_26_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1583) | ~rob_val_1_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1039)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_26_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_26_br_mask <= rob_uop_1_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1040) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_27_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_27_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_27_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_27_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_27_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_27_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_27_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_27_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_27_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_27_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_27_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_27_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_27_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_27_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_27_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_27_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1584) | ~rob_val_1_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1040)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_27_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_27_br_mask <= rob_uop_1_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1041) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_28_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_28_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_28_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_28_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_28_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_28_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_28_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_28_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_28_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_28_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_28_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_28_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_28_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_28_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_28_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_28_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1585) | ~rob_val_1_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1041)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_28_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_28_br_mask <= rob_uop_1_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1042) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_29_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_29_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_29_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_29_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_29_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_29_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_29_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_29_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_29_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_29_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_29_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_29_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_29_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_29_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_29_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_29_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1586) | ~rob_val_1_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1042)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_29_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_29_br_mask <= rob_uop_1_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1043) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_30_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_30_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_30_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_30_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_30_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_30_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_30_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_30_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_30_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_30_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_30_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_30_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_30_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_30_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_30_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_30_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1587) | ~rob_val_1_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1043)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_30_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_30_br_mask <= rob_uop_1_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1044) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_1_31_uopc <= io_enq_uops_1_uopc;	// rob.scala:310:28
      rob_uop_1_31_is_rvc <= io_enq_uops_1_is_rvc;	// rob.scala:310:28
      rob_uop_1_31_ftq_idx <= io_enq_uops_1_ftq_idx;	// rob.scala:310:28
      rob_uop_1_31_edge_inst <= io_enq_uops_1_edge_inst;	// rob.scala:310:28
      rob_uop_1_31_pc_lob <= io_enq_uops_1_pc_lob;	// rob.scala:310:28
      rob_uop_1_31_pdst <= io_enq_uops_1_pdst;	// rob.scala:310:28
      rob_uop_1_31_stale_pdst <= io_enq_uops_1_stale_pdst;	// rob.scala:310:28
      rob_uop_1_31_is_fencei <= io_enq_uops_1_is_fencei;	// rob.scala:310:28
      rob_uop_1_31_uses_ldq <= io_enq_uops_1_uses_ldq;	// rob.scala:310:28
      rob_uop_1_31_uses_stq <= io_enq_uops_1_uses_stq;	// rob.scala:310:28
      rob_uop_1_31_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_1_31_flush_on_commit <= io_enq_uops_1_flush_on_commit;	// rob.scala:310:28
      rob_uop_1_31_ldst <= io_enq_uops_1_ldst;	// rob.scala:310:28
      rob_uop_1_31_ldst_val <= io_enq_uops_1_ldst_val;	// rob.scala:310:28
      rob_uop_1_31_dst_rtype <= io_enq_uops_1_dst_rtype;	// rob.scala:310:28
      rob_uop_1_31_fp_val <= io_enq_uops_1_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_1588) | ~rob_val_1_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1044)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_1_31_br_mask <= io_enq_uops_1_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_1_31_br_mask <= rob_uop_1_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_1_0 <=
      ~_GEN_1525
      & (_GEN_39 & _GEN_887 | (_GEN_1013 ? io_enq_uops_1_exception : rob_exception_1_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_1 <=
      ~_GEN_1526
      & (_GEN_39 & _GEN_888 | (_GEN_1014 ? io_enq_uops_1_exception : rob_exception_1_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_2 <=
      ~_GEN_1527
      & (_GEN_39 & _GEN_889 | (_GEN_1015 ? io_enq_uops_1_exception : rob_exception_1_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_3 <=
      ~_GEN_1528
      & (_GEN_39 & _GEN_890 | (_GEN_1016 ? io_enq_uops_1_exception : rob_exception_1_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_4 <=
      ~_GEN_1529
      & (_GEN_39 & _GEN_891 | (_GEN_1017 ? io_enq_uops_1_exception : rob_exception_1_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_5 <=
      ~_GEN_1530
      & (_GEN_39 & _GEN_892 | (_GEN_1018 ? io_enq_uops_1_exception : rob_exception_1_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_6 <=
      ~_GEN_1531
      & (_GEN_39 & _GEN_893 | (_GEN_1019 ? io_enq_uops_1_exception : rob_exception_1_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_7 <=
      ~_GEN_1532
      & (_GEN_39 & _GEN_894 | (_GEN_1020 ? io_enq_uops_1_exception : rob_exception_1_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_8 <=
      ~_GEN_1533
      & (_GEN_39 & _GEN_895 | (_GEN_1021 ? io_enq_uops_1_exception : rob_exception_1_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_9 <=
      ~_GEN_1534
      & (_GEN_39 & _GEN_896 | (_GEN_1022 ? io_enq_uops_1_exception : rob_exception_1_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_10 <=
      ~_GEN_1535
      & (_GEN_39 & _GEN_897 | (_GEN_1023 ? io_enq_uops_1_exception : rob_exception_1_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_11 <=
      ~_GEN_1536
      & (_GEN_39 & _GEN_898 | (_GEN_1024 ? io_enq_uops_1_exception : rob_exception_1_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_12 <=
      ~_GEN_1537
      & (_GEN_39 & _GEN_899 | (_GEN_1025 ? io_enq_uops_1_exception : rob_exception_1_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_13 <=
      ~_GEN_1538
      & (_GEN_39 & _GEN_900 | (_GEN_1026 ? io_enq_uops_1_exception : rob_exception_1_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_14 <=
      ~_GEN_1539
      & (_GEN_39 & _GEN_901 | (_GEN_1027 ? io_enq_uops_1_exception : rob_exception_1_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_15 <=
      ~_GEN_1540
      & (_GEN_39 & _GEN_902 | (_GEN_1028 ? io_enq_uops_1_exception : rob_exception_1_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_16 <=
      ~_GEN_1541
      & (_GEN_39 & _GEN_903 | (_GEN_1029 ? io_enq_uops_1_exception : rob_exception_1_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_17 <=
      ~_GEN_1542
      & (_GEN_39 & _GEN_904 | (_GEN_1030 ? io_enq_uops_1_exception : rob_exception_1_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_18 <=
      ~_GEN_1543
      & (_GEN_39 & _GEN_905 | (_GEN_1031 ? io_enq_uops_1_exception : rob_exception_1_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_19 <=
      ~_GEN_1544
      & (_GEN_39 & _GEN_906 | (_GEN_1032 ? io_enq_uops_1_exception : rob_exception_1_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_20 <=
      ~_GEN_1545
      & (_GEN_39 & _GEN_907 | (_GEN_1033 ? io_enq_uops_1_exception : rob_exception_1_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_21 <=
      ~_GEN_1546
      & (_GEN_39 & _GEN_908 | (_GEN_1034 ? io_enq_uops_1_exception : rob_exception_1_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_22 <=
      ~_GEN_1547
      & (_GEN_39 & _GEN_909 | (_GEN_1035 ? io_enq_uops_1_exception : rob_exception_1_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_23 <=
      ~_GEN_1548
      & (_GEN_39 & _GEN_910 | (_GEN_1036 ? io_enq_uops_1_exception : rob_exception_1_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_24 <=
      ~_GEN_1549
      & (_GEN_39 & _GEN_911 | (_GEN_1037 ? io_enq_uops_1_exception : rob_exception_1_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_25 <=
      ~_GEN_1550
      & (_GEN_39 & _GEN_912 | (_GEN_1038 ? io_enq_uops_1_exception : rob_exception_1_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_26 <=
      ~_GEN_1551
      & (_GEN_39 & _GEN_913 | (_GEN_1039 ? io_enq_uops_1_exception : rob_exception_1_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_27 <=
      ~_GEN_1552
      & (_GEN_39 & _GEN_914 | (_GEN_1040 ? io_enq_uops_1_exception : rob_exception_1_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_28 <=
      ~_GEN_1553
      & (_GEN_39 & _GEN_915 | (_GEN_1041 ? io_enq_uops_1_exception : rob_exception_1_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_29 <=
      ~_GEN_1554
      & (_GEN_39 & _GEN_916 | (_GEN_1042 ? io_enq_uops_1_exception : rob_exception_1_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_30 <=
      ~_GEN_1555
      & (_GEN_39 & _GEN_917 | (_GEN_1043 ? io_enq_uops_1_exception : rob_exception_1_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_1_31 <=
      ~_GEN_1556
      & (_GEN_39 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_1044 ? io_enq_uops_1_exception : rob_exception_1_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_1_0 <=
      ~(_GEN_35 & _GEN_666)
      & (_GEN_1365
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_476 | _GEN_1237 | _GEN_31 & _GEN_286)
             & (_GEN_1109
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1013 & rob_predicated_1_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_1 <=
      ~(_GEN_35 & _GEN_669)
      & (_GEN_1366
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_479 | _GEN_1238 | _GEN_31 & _GEN_289)
             & (_GEN_1110
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1014 & rob_predicated_1_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_2 <=
      ~(_GEN_35 & _GEN_672)
      & (_GEN_1367
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_482 | _GEN_1239 | _GEN_31 & _GEN_292)
             & (_GEN_1111
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1015 & rob_predicated_1_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_3 <=
      ~(_GEN_35 & _GEN_675)
      & (_GEN_1368
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_485 | _GEN_1240 | _GEN_31 & _GEN_295)
             & (_GEN_1112
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1016 & rob_predicated_1_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_4 <=
      ~(_GEN_35 & _GEN_678)
      & (_GEN_1369
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_488 | _GEN_1241 | _GEN_31 & _GEN_298)
             & (_GEN_1113
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1017 & rob_predicated_1_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_5 <=
      ~(_GEN_35 & _GEN_681)
      & (_GEN_1370
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_491 | _GEN_1242 | _GEN_31 & _GEN_301)
             & (_GEN_1114
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1018 & rob_predicated_1_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_6 <=
      ~(_GEN_35 & _GEN_684)
      & (_GEN_1371
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_494 | _GEN_1243 | _GEN_31 & _GEN_304)
             & (_GEN_1115
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1019 & rob_predicated_1_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_7 <=
      ~(_GEN_35 & _GEN_687)
      & (_GEN_1372
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_497 | _GEN_1244 | _GEN_31 & _GEN_307)
             & (_GEN_1116
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1020 & rob_predicated_1_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_8 <=
      ~(_GEN_35 & _GEN_690)
      & (_GEN_1373
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_500 | _GEN_1245 | _GEN_31 & _GEN_310)
             & (_GEN_1117
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1021 & rob_predicated_1_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_9 <=
      ~(_GEN_35 & _GEN_693)
      & (_GEN_1374
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_503 | _GEN_1246 | _GEN_31 & _GEN_313)
             & (_GEN_1118
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1022 & rob_predicated_1_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_10 <=
      ~(_GEN_35 & _GEN_696)
      & (_GEN_1375
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_506 | _GEN_1247 | _GEN_31 & _GEN_316)
             & (_GEN_1119
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1023 & rob_predicated_1_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_11 <=
      ~(_GEN_35 & _GEN_699)
      & (_GEN_1376
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_509 | _GEN_1248 | _GEN_31 & _GEN_319)
             & (_GEN_1120
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1024 & rob_predicated_1_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_12 <=
      ~(_GEN_35 & _GEN_702)
      & (_GEN_1377
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_512 | _GEN_1249 | _GEN_31 & _GEN_322)
             & (_GEN_1121
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1025 & rob_predicated_1_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_13 <=
      ~(_GEN_35 & _GEN_705)
      & (_GEN_1378
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_515 | _GEN_1250 | _GEN_31 & _GEN_325)
             & (_GEN_1122
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1026 & rob_predicated_1_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_14 <=
      ~(_GEN_35 & _GEN_708)
      & (_GEN_1379
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_518 | _GEN_1251 | _GEN_31 & _GEN_328)
             & (_GEN_1123
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1027 & rob_predicated_1_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_15 <=
      ~(_GEN_35 & _GEN_711)
      & (_GEN_1380
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_521 | _GEN_1252 | _GEN_31 & _GEN_331)
             & (_GEN_1124
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1028 & rob_predicated_1_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_16 <=
      ~(_GEN_35 & _GEN_714)
      & (_GEN_1381
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_524 | _GEN_1253 | _GEN_31 & _GEN_334)
             & (_GEN_1125
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1029 & rob_predicated_1_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_17 <=
      ~(_GEN_35 & _GEN_717)
      & (_GEN_1382
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_527 | _GEN_1254 | _GEN_31 & _GEN_337)
             & (_GEN_1126
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1030 & rob_predicated_1_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_18 <=
      ~(_GEN_35 & _GEN_720)
      & (_GEN_1383
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_530 | _GEN_1255 | _GEN_31 & _GEN_340)
             & (_GEN_1127
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1031 & rob_predicated_1_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_19 <=
      ~(_GEN_35 & _GEN_723)
      & (_GEN_1384
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_533 | _GEN_1256 | _GEN_31 & _GEN_343)
             & (_GEN_1128
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1032 & rob_predicated_1_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_20 <=
      ~(_GEN_35 & _GEN_726)
      & (_GEN_1385
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_536 | _GEN_1257 | _GEN_31 & _GEN_346)
             & (_GEN_1129
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1033 & rob_predicated_1_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_21 <=
      ~(_GEN_35 & _GEN_729)
      & (_GEN_1386
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_539 | _GEN_1258 | _GEN_31 & _GEN_349)
             & (_GEN_1130
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1034 & rob_predicated_1_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_22 <=
      ~(_GEN_35 & _GEN_732)
      & (_GEN_1387
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_542 | _GEN_1259 | _GEN_31 & _GEN_352)
             & (_GEN_1131
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1035 & rob_predicated_1_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_23 <=
      ~(_GEN_35 & _GEN_735)
      & (_GEN_1388
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_545 | _GEN_1260 | _GEN_31 & _GEN_355)
             & (_GEN_1132
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1036 & rob_predicated_1_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_24 <=
      ~(_GEN_35 & _GEN_738)
      & (_GEN_1389
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_548 | _GEN_1261 | _GEN_31 & _GEN_358)
             & (_GEN_1133
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1037 & rob_predicated_1_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_25 <=
      ~(_GEN_35 & _GEN_741)
      & (_GEN_1390
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_551 | _GEN_1262 | _GEN_31 & _GEN_361)
             & (_GEN_1134
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1038 & rob_predicated_1_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_26 <=
      ~(_GEN_35 & _GEN_744)
      & (_GEN_1391
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_554 | _GEN_1263 | _GEN_31 & _GEN_364)
             & (_GEN_1135
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1039 & rob_predicated_1_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_27 <=
      ~(_GEN_35 & _GEN_747)
      & (_GEN_1392
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_557 | _GEN_1264 | _GEN_31 & _GEN_367)
             & (_GEN_1136
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1040 & rob_predicated_1_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_28 <=
      ~(_GEN_35 & _GEN_750)
      & (_GEN_1393
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_560 | _GEN_1265 | _GEN_31 & _GEN_370)
             & (_GEN_1137
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1041 & rob_predicated_1_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_29 <=
      ~(_GEN_35 & _GEN_753)
      & (_GEN_1394
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_563 | _GEN_1266 | _GEN_31 & _GEN_373)
             & (_GEN_1138
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1042 & rob_predicated_1_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_30 <=
      ~(_GEN_35 & _GEN_756)
      & (_GEN_1395
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & _GEN_566 | _GEN_1267 | _GEN_31 & _GEN_376)
             & (_GEN_1139
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1043 & rob_predicated_1_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_1_31 <=
      ~(_GEN_35 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])))
      & (_GEN_1396
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_33 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1268 | _GEN_31
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_1140
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1044 & rob_predicated_1_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    if (_GEN_68) begin	// rob.scala:361:31
      automatic logic _GEN_2467;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2468;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2469;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2470;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2471;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2472;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2473;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2474;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2475;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2476;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2477;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2478;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2479;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2480;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2481;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2482;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2483;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2484;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2485;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2486;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2487;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2488;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2489;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2490;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2491;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2492;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2493;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2494;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2495;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2496;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2497;	// rob.scala:346:69, :361:75, :363:26
      automatic logic _GEN_2498;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2467 = _GEN_856 | _GEN_2069;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2468 = _GEN_857 | _GEN_2070;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2469 = _GEN_858 | _GEN_2071;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2470 = _GEN_859 | _GEN_2072;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2471 = _GEN_860 | _GEN_2073;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2472 = _GEN_861 | _GEN_2074;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2473 = _GEN_862 | _GEN_2075;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2474 = _GEN_863 | _GEN_2076;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2475 = _GEN_864 | _GEN_2077;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2476 = _GEN_865 | _GEN_2078;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2477 = _GEN_866 | _GEN_2079;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2478 = _GEN_867 | _GEN_2080;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2479 = _GEN_868 | _GEN_2081;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2480 = _GEN_869 | _GEN_2082;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2481 = _GEN_870 | _GEN_2083;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2482 = _GEN_871 | _GEN_2084;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2483 = _GEN_872 | _GEN_2085;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2484 = _GEN_873 | _GEN_2086;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2485 = _GEN_874 | _GEN_2087;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2486 = _GEN_875 | _GEN_2088;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2487 = _GEN_876 | _GEN_2089;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2488 = _GEN_877 | _GEN_2090;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2489 = _GEN_878 | _GEN_2091;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2490 = _GEN_879 | _GEN_2092;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2491 = _GEN_880 | _GEN_2093;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2492 = _GEN_881 | _GEN_2094;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2493 = _GEN_882 | _GEN_2095;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2494 = _GEN_883 | _GEN_2096;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2495 = _GEN_884 | _GEN_2097;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2496 = _GEN_885 | _GEN_2098;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2497 = _GEN_886 | _GEN_2099;	// rob.scala:346:69, :361:75, :363:26
      _GEN_2498 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_2100;	// rob.scala:236:31, :268:25, :346:69, :361:75, :363:26
      rob_bsy_2_0 <= ~_GEN_2467 & _GEN_1974;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_1 <= ~_GEN_2468 & _GEN_1976;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_2 <= ~_GEN_2469 & _GEN_1978;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_3 <= ~_GEN_2470 & _GEN_1980;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_4 <= ~_GEN_2471 & _GEN_1982;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_5 <= ~_GEN_2472 & _GEN_1984;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_6 <= ~_GEN_2473 & _GEN_1986;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_7 <= ~_GEN_2474 & _GEN_1988;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_8 <= ~_GEN_2475 & _GEN_1990;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_9 <= ~_GEN_2476 & _GEN_1992;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_10 <= ~_GEN_2477 & _GEN_1994;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_11 <= ~_GEN_2478 & _GEN_1996;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_12 <= ~_GEN_2479 & _GEN_1998;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_13 <= ~_GEN_2480 & _GEN_2000;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_14 <= ~_GEN_2481 & _GEN_2002;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_15 <= ~_GEN_2482 & _GEN_2004;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_16 <= ~_GEN_2483 & _GEN_2006;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_17 <= ~_GEN_2484 & _GEN_2008;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_18 <= ~_GEN_2485 & _GEN_2010;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_19 <= ~_GEN_2486 & _GEN_2012;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_20 <= ~_GEN_2487 & _GEN_2014;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_21 <= ~_GEN_2488 & _GEN_2016;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_22 <= ~_GEN_2489 & _GEN_2018;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_23 <= ~_GEN_2490 & _GEN_2020;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_24 <= ~_GEN_2491 & _GEN_2022;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_25 <= ~_GEN_2492 & _GEN_2024;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_26 <= ~_GEN_2493 & _GEN_2026;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_27 <= ~_GEN_2494 & _GEN_2028;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_28 <= ~_GEN_2495 & _GEN_2030;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_29 <= ~_GEN_2496 & _GEN_2032;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_30 <= ~_GEN_2497 & _GEN_2034;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_31 <= ~_GEN_2498 & _GEN_2036;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_unsafe_2_0 <= ~_GEN_2467 & _GEN_2037;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_1 <= ~_GEN_2468 & _GEN_2038;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_2 <= ~_GEN_2469 & _GEN_2039;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_3 <= ~_GEN_2470 & _GEN_2040;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_4 <= ~_GEN_2471 & _GEN_2041;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_5 <= ~_GEN_2472 & _GEN_2042;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_6 <= ~_GEN_2473 & _GEN_2043;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_7 <= ~_GEN_2474 & _GEN_2044;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_8 <= ~_GEN_2475 & _GEN_2045;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_9 <= ~_GEN_2476 & _GEN_2046;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_10 <= ~_GEN_2477 & _GEN_2047;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_11 <= ~_GEN_2478 & _GEN_2048;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_12 <= ~_GEN_2479 & _GEN_2049;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_13 <= ~_GEN_2480 & _GEN_2050;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_14 <= ~_GEN_2481 & _GEN_2051;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_15 <= ~_GEN_2482 & _GEN_2052;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_16 <= ~_GEN_2483 & _GEN_2053;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_17 <= ~_GEN_2484 & _GEN_2054;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_18 <= ~_GEN_2485 & _GEN_2055;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_19 <= ~_GEN_2486 & _GEN_2056;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_20 <= ~_GEN_2487 & _GEN_2057;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_21 <= ~_GEN_2488 & _GEN_2058;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_22 <= ~_GEN_2489 & _GEN_2059;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_23 <= ~_GEN_2490 & _GEN_2060;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_24 <= ~_GEN_2491 & _GEN_2061;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_25 <= ~_GEN_2492 & _GEN_2062;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_26 <= ~_GEN_2493 & _GEN_2063;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_27 <= ~_GEN_2494 & _GEN_2064;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_28 <= ~_GEN_2495 & _GEN_2065;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_29 <= ~_GEN_2496 & _GEN_2066;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_30 <= ~_GEN_2497 & _GEN_2067;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_31 <= ~_GEN_2498 & _GEN_2068;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
    end
    else begin	// rob.scala:361:31
      rob_bsy_2_0 <= ~_GEN_2069 & _GEN_1974;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_1 <= ~_GEN_2070 & _GEN_1976;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_2 <= ~_GEN_2071 & _GEN_1978;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_3 <= ~_GEN_2072 & _GEN_1980;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_4 <= ~_GEN_2073 & _GEN_1982;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_5 <= ~_GEN_2074 & _GEN_1984;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_6 <= ~_GEN_2075 & _GEN_1986;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_7 <= ~_GEN_2076 & _GEN_1988;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_8 <= ~_GEN_2077 & _GEN_1990;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_9 <= ~_GEN_2078 & _GEN_1992;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_10 <= ~_GEN_2079 & _GEN_1994;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_11 <= ~_GEN_2080 & _GEN_1996;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_12 <= ~_GEN_2081 & _GEN_1998;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_13 <= ~_GEN_2082 & _GEN_2000;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_14 <= ~_GEN_2083 & _GEN_2002;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_15 <= ~_GEN_2084 & _GEN_2004;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_16 <= ~_GEN_2085 & _GEN_2006;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_17 <= ~_GEN_2086 & _GEN_2008;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_18 <= ~_GEN_2087 & _GEN_2010;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_19 <= ~_GEN_2088 & _GEN_2012;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_20 <= ~_GEN_2089 & _GEN_2014;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_21 <= ~_GEN_2090 & _GEN_2016;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_22 <= ~_GEN_2091 & _GEN_2018;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_23 <= ~_GEN_2092 & _GEN_2020;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_24 <= ~_GEN_2093 & _GEN_2022;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_25 <= ~_GEN_2094 & _GEN_2024;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_26 <= ~_GEN_2095 & _GEN_2026;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_27 <= ~_GEN_2096 & _GEN_2028;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_28 <= ~_GEN_2097 & _GEN_2030;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_29 <= ~_GEN_2098 & _GEN_2032;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_30 <= ~_GEN_2099 & _GEN_2034;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_bsy_2_31 <= ~_GEN_2100 & _GEN_2036;	// rob.scala:308:28, :346:69, :347:31, :361:75, :363:26
      rob_unsafe_2_0 <= ~_GEN_2069 & _GEN_2037;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_1 <= ~_GEN_2070 & _GEN_2038;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_2 <= ~_GEN_2071 & _GEN_2039;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_3 <= ~_GEN_2072 & _GEN_2040;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_4 <= ~_GEN_2073 & _GEN_2041;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_5 <= ~_GEN_2074 & _GEN_2042;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_6 <= ~_GEN_2075 & _GEN_2043;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_7 <= ~_GEN_2076 & _GEN_2044;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_8 <= ~_GEN_2077 & _GEN_2045;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_9 <= ~_GEN_2078 & _GEN_2046;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_10 <= ~_GEN_2079 & _GEN_2047;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_11 <= ~_GEN_2080 & _GEN_2048;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_12 <= ~_GEN_2081 & _GEN_2049;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_13 <= ~_GEN_2082 & _GEN_2050;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_14 <= ~_GEN_2083 & _GEN_2051;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_15 <= ~_GEN_2084 & _GEN_2052;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_16 <= ~_GEN_2085 & _GEN_2053;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_17 <= ~_GEN_2086 & _GEN_2054;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_18 <= ~_GEN_2087 & _GEN_2055;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_19 <= ~_GEN_2088 & _GEN_2056;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_20 <= ~_GEN_2089 & _GEN_2057;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_21 <= ~_GEN_2090 & _GEN_2058;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_22 <= ~_GEN_2091 & _GEN_2059;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_23 <= ~_GEN_2092 & _GEN_2060;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_24 <= ~_GEN_2093 & _GEN_2061;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_25 <= ~_GEN_2094 & _GEN_2062;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_26 <= ~_GEN_2095 & _GEN_2063;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_27 <= ~_GEN_2096 & _GEN_2064;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_28 <= ~_GEN_2097 & _GEN_2065;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_29 <= ~_GEN_2098 & _GEN_2066;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_30 <= ~_GEN_2099 & _GEN_2067;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
      rob_unsafe_2_31 <= ~_GEN_2100 & _GEN_2068;	// rob.scala:309:28, :346:69, :348:31, :361:75, :363:26, :364:26
    end
    if (_GEN_1589) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_0_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_0_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_0_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_0_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_0_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_0_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_0_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_0_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_0_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_0_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_0_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_0_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_0_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_0_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_0_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_0_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2133) | ~rob_val_2_0) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1589)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_0_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_0_br_mask <= rob_uop_2_0_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1590) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_1_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_1_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_1_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_1_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_1_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_1_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_1_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_1_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_1_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_1_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_1_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_1_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_1_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_1_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_1_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_1_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2134) | ~rob_val_2_1) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1590)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_1_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_1_br_mask <= rob_uop_2_1_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1591) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_2_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_2_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_2_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_2_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_2_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_2_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_2_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_2_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_2_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_2_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_2_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_2_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_2_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_2_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_2_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_2_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2135) | ~rob_val_2_2) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1591)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_2_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_2_br_mask <= rob_uop_2_2_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1592) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_3_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_3_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_3_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_3_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_3_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_3_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_3_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_3_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_3_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_3_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_3_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_3_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_3_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_3_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_3_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_3_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2136) | ~rob_val_2_3) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1592)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_3_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_3_br_mask <= rob_uop_2_3_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1593) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_4_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_4_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_4_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_4_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_4_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_4_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_4_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_4_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_4_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_4_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_4_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_4_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_4_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_4_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_4_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_4_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2137) | ~rob_val_2_4) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1593)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_4_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_4_br_mask <= rob_uop_2_4_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1594) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_5_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_5_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_5_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_5_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_5_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_5_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_5_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_5_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_5_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_5_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_5_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_5_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_5_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_5_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_5_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_5_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2138) | ~rob_val_2_5) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1594)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_5_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_5_br_mask <= rob_uop_2_5_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1595) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_6_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_6_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_6_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_6_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_6_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_6_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_6_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_6_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_6_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_6_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_6_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_6_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_6_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_6_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_6_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_6_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2139) | ~rob_val_2_6) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1595)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_6_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_6_br_mask <= rob_uop_2_6_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1596) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_7_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_7_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_7_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_7_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_7_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_7_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_7_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_7_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_7_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_7_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_7_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_7_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_7_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_7_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_7_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_7_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2140) | ~rob_val_2_7) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1596)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_7_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_7_br_mask <= rob_uop_2_7_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1597) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_8_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_8_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_8_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_8_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_8_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_8_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_8_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_8_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_8_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_8_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_8_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_8_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_8_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_8_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_8_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_8_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2141) | ~rob_val_2_8) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1597)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_8_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_8_br_mask <= rob_uop_2_8_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1598) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_9_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_9_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_9_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_9_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_9_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_9_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_9_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_9_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_9_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_9_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_9_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_9_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_9_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_9_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_9_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_9_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2142) | ~rob_val_2_9) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1598)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_9_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_9_br_mask <= rob_uop_2_9_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1599) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_10_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_10_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_10_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_10_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_10_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_10_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_10_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_10_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_10_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_10_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_10_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_10_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_10_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_10_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_10_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_10_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2143) | ~rob_val_2_10) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1599)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_10_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_10_br_mask <= rob_uop_2_10_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1600) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_11_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_11_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_11_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_11_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_11_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_11_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_11_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_11_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_11_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_11_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_11_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_11_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_11_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_11_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_11_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_11_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2144) | ~rob_val_2_11) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1600)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_11_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_11_br_mask <= rob_uop_2_11_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1601) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_12_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_12_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_12_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_12_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_12_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_12_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_12_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_12_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_12_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_12_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_12_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_12_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_12_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_12_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_12_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_12_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2145) | ~rob_val_2_12) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1601)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_12_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_12_br_mask <= rob_uop_2_12_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1602) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_13_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_13_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_13_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_13_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_13_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_13_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_13_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_13_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_13_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_13_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_13_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_13_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_13_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_13_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_13_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_13_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2146) | ~rob_val_2_13) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1602)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_13_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_13_br_mask <= rob_uop_2_13_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1603) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_14_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_14_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_14_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_14_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_14_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_14_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_14_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_14_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_14_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_14_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_14_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_14_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_14_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_14_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_14_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_14_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2147) | ~rob_val_2_14) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1603)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_14_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_14_br_mask <= rob_uop_2_14_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1604) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_15_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_15_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_15_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_15_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_15_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_15_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_15_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_15_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_15_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_15_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_15_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_15_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_15_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_15_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_15_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_15_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2148) | ~rob_val_2_15) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1604)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_15_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_15_br_mask <= rob_uop_2_15_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1605) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_16_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_16_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_16_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_16_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_16_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_16_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_16_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_16_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_16_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_16_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_16_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_16_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_16_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_16_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_16_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_16_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2149) | ~rob_val_2_16) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1605)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_16_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_16_br_mask <= rob_uop_2_16_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1606) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_17_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_17_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_17_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_17_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_17_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_17_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_17_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_17_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_17_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_17_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_17_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_17_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_17_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_17_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_17_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_17_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2150) | ~rob_val_2_17) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1606)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_17_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_17_br_mask <= rob_uop_2_17_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1607) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_18_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_18_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_18_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_18_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_18_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_18_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_18_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_18_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_18_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_18_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_18_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_18_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_18_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_18_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_18_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_18_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2151) | ~rob_val_2_18) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1607)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_18_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_18_br_mask <= rob_uop_2_18_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1608) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_19_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_19_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_19_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_19_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_19_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_19_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_19_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_19_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_19_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_19_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_19_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_19_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_19_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_19_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_19_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_19_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2152) | ~rob_val_2_19) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1608)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_19_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_19_br_mask <= rob_uop_2_19_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1609) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_20_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_20_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_20_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_20_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_20_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_20_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_20_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_20_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_20_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_20_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_20_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_20_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_20_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_20_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_20_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_20_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2153) | ~rob_val_2_20) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1609)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_20_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_20_br_mask <= rob_uop_2_20_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1610) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_21_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_21_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_21_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_21_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_21_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_21_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_21_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_21_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_21_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_21_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_21_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_21_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_21_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_21_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_21_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_21_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2154) | ~rob_val_2_21) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1610)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_21_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_21_br_mask <= rob_uop_2_21_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1611) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_22_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_22_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_22_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_22_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_22_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_22_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_22_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_22_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_22_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_22_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_22_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_22_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_22_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_22_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_22_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_22_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2155) | ~rob_val_2_22) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1611)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_22_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_22_br_mask <= rob_uop_2_22_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1612) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_23_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_23_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_23_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_23_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_23_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_23_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_23_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_23_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_23_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_23_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_23_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_23_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_23_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_23_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_23_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_23_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2156) | ~rob_val_2_23) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1612)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_23_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_23_br_mask <= rob_uop_2_23_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1613) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_24_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_24_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_24_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_24_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_24_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_24_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_24_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_24_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_24_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_24_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_24_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_24_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_24_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_24_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_24_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_24_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2157) | ~rob_val_2_24) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1613)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_24_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_24_br_mask <= rob_uop_2_24_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1614) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_25_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_25_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_25_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_25_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_25_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_25_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_25_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_25_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_25_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_25_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_25_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_25_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_25_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_25_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_25_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_25_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2158) | ~rob_val_2_25) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1614)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_25_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_25_br_mask <= rob_uop_2_25_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1615) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_26_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_26_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_26_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_26_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_26_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_26_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_26_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_26_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_26_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_26_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_26_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_26_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_26_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_26_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_26_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_26_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2159) | ~rob_val_2_26) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1615)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_26_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_26_br_mask <= rob_uop_2_26_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1616) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_27_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_27_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_27_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_27_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_27_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_27_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_27_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_27_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_27_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_27_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_27_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_27_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_27_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_27_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_27_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_27_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2160) | ~rob_val_2_27) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1616)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_27_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_27_br_mask <= rob_uop_2_27_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1617) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_28_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_28_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_28_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_28_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_28_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_28_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_28_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_28_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_28_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_28_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_28_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_28_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_28_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_28_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_28_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_28_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2161) | ~rob_val_2_28) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1617)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_28_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_28_br_mask <= rob_uop_2_28_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1618) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_29_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_29_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_29_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_29_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_29_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_29_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_29_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_29_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_29_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_29_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_29_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_29_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_29_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_29_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_29_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_29_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2162) | ~rob_val_2_29) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1618)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_29_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_29_br_mask <= rob_uop_2_29_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1619) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_30_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_30_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_30_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_30_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_30_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_30_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_30_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_30_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_30_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_30_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_30_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_30_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_30_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_30_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_30_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_30_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2163) | ~rob_val_2_30) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1619)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_30_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_30_br_mask <= rob_uop_2_30_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    if (_GEN_1620) begin	// rob.scala:307:32, :323:29, :324:31
      rob_uop_2_31_uopc <= io_enq_uops_2_uopc;	// rob.scala:310:28
      rob_uop_2_31_is_rvc <= io_enq_uops_2_is_rvc;	// rob.scala:310:28
      rob_uop_2_31_ftq_idx <= io_enq_uops_2_ftq_idx;	// rob.scala:310:28
      rob_uop_2_31_edge_inst <= io_enq_uops_2_edge_inst;	// rob.scala:310:28
      rob_uop_2_31_pc_lob <= io_enq_uops_2_pc_lob;	// rob.scala:310:28
      rob_uop_2_31_pdst <= io_enq_uops_2_pdst;	// rob.scala:310:28
      rob_uop_2_31_stale_pdst <= io_enq_uops_2_stale_pdst;	// rob.scala:310:28
      rob_uop_2_31_is_fencei <= io_enq_uops_2_is_fencei;	// rob.scala:310:28
      rob_uop_2_31_uses_ldq <= io_enq_uops_2_uses_ldq;	// rob.scala:310:28
      rob_uop_2_31_uses_stq <= io_enq_uops_2_uses_stq;	// rob.scala:310:28
      rob_uop_2_31_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;	// rob.scala:310:28
      rob_uop_2_31_flush_on_commit <= io_enq_uops_2_flush_on_commit;	// rob.scala:310:28
      rob_uop_2_31_ldst <= io_enq_uops_2_ldst;	// rob.scala:310:28
      rob_uop_2_31_ldst_val <= io_enq_uops_2_ldst_val;	// rob.scala:310:28
      rob_uop_2_31_dst_rtype <= io_enq_uops_2_dst_rtype;	// rob.scala:310:28
      rob_uop_2_31_fp_val <= io_enq_uops_2_fp_val;	// rob.scala:310:28
    end
    if ((|_GEN_2164) | ~rob_val_2_31) begin	// rob.scala:307:32, :323:29, :455:7, :458:32, util.scala:118:{51,59}
      if (_GEN_1620)	// rob.scala:307:32, :323:29, :324:31
        rob_uop_2_31_br_mask <= io_enq_uops_2_br_mask;	// rob.scala:310:28
    end
    else	// rob.scala:323:29, :455:7, :458:32
      rob_uop_2_31_br_mask <= rob_uop_2_31_br_mask & ~io_brupdate_b1_resolve_mask;	// rob.scala:310:28, util.scala:89:{21,23}
    rob_exception_2_0 <=
      ~_GEN_2101
      & (_GEN_69 & _GEN_887 | (_GEN_1589 ? io_enq_uops_2_exception : rob_exception_2_0));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_1 <=
      ~_GEN_2102
      & (_GEN_69 & _GEN_888 | (_GEN_1590 ? io_enq_uops_2_exception : rob_exception_2_1));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_2 <=
      ~_GEN_2103
      & (_GEN_69 & _GEN_889 | (_GEN_1591 ? io_enq_uops_2_exception : rob_exception_2_2));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_3 <=
      ~_GEN_2104
      & (_GEN_69 & _GEN_890 | (_GEN_1592 ? io_enq_uops_2_exception : rob_exception_2_3));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_4 <=
      ~_GEN_2105
      & (_GEN_69 & _GEN_891 | (_GEN_1593 ? io_enq_uops_2_exception : rob_exception_2_4));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_5 <=
      ~_GEN_2106
      & (_GEN_69 & _GEN_892 | (_GEN_1594 ? io_enq_uops_2_exception : rob_exception_2_5));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_6 <=
      ~_GEN_2107
      & (_GEN_69 & _GEN_893 | (_GEN_1595 ? io_enq_uops_2_exception : rob_exception_2_6));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_7 <=
      ~_GEN_2108
      & (_GEN_69 & _GEN_894 | (_GEN_1596 ? io_enq_uops_2_exception : rob_exception_2_7));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_8 <=
      ~_GEN_2109
      & (_GEN_69 & _GEN_895 | (_GEN_1597 ? io_enq_uops_2_exception : rob_exception_2_8));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_9 <=
      ~_GEN_2110
      & (_GEN_69 & _GEN_896 | (_GEN_1598 ? io_enq_uops_2_exception : rob_exception_2_9));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_10 <=
      ~_GEN_2111
      & (_GEN_69 & _GEN_897 | (_GEN_1599 ? io_enq_uops_2_exception : rob_exception_2_10));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_11 <=
      ~_GEN_2112
      & (_GEN_69 & _GEN_898 | (_GEN_1600 ? io_enq_uops_2_exception : rob_exception_2_11));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_12 <=
      ~_GEN_2113
      & (_GEN_69 & _GEN_899 | (_GEN_1601 ? io_enq_uops_2_exception : rob_exception_2_12));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_13 <=
      ~_GEN_2114
      & (_GEN_69 & _GEN_900 | (_GEN_1602 ? io_enq_uops_2_exception : rob_exception_2_13));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_14 <=
      ~_GEN_2115
      & (_GEN_69 & _GEN_901 | (_GEN_1603 ? io_enq_uops_2_exception : rob_exception_2_14));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_15 <=
      ~_GEN_2116
      & (_GEN_69 & _GEN_902 | (_GEN_1604 ? io_enq_uops_2_exception : rob_exception_2_15));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_16 <=
      ~_GEN_2117
      & (_GEN_69 & _GEN_903 | (_GEN_1605 ? io_enq_uops_2_exception : rob_exception_2_16));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_17 <=
      ~_GEN_2118
      & (_GEN_69 & _GEN_904 | (_GEN_1606 ? io_enq_uops_2_exception : rob_exception_2_17));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_18 <=
      ~_GEN_2119
      & (_GEN_69 & _GEN_905 | (_GEN_1607 ? io_enq_uops_2_exception : rob_exception_2_18));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_19 <=
      ~_GEN_2120
      & (_GEN_69 & _GEN_906 | (_GEN_1608 ? io_enq_uops_2_exception : rob_exception_2_19));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_20 <=
      ~_GEN_2121
      & (_GEN_69 & _GEN_907 | (_GEN_1609 ? io_enq_uops_2_exception : rob_exception_2_20));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_21 <=
      ~_GEN_2122
      & (_GEN_69 & _GEN_908 | (_GEN_1610 ? io_enq_uops_2_exception : rob_exception_2_21));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_22 <=
      ~_GEN_2123
      & (_GEN_69 & _GEN_909 | (_GEN_1611 ? io_enq_uops_2_exception : rob_exception_2_22));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_23 <=
      ~_GEN_2124
      & (_GEN_69 & _GEN_910 | (_GEN_1612 ? io_enq_uops_2_exception : rob_exception_2_23));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_24 <=
      ~_GEN_2125
      & (_GEN_69 & _GEN_911 | (_GEN_1613 ? io_enq_uops_2_exception : rob_exception_2_24));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_25 <=
      ~_GEN_2126
      & (_GEN_69 & _GEN_912 | (_GEN_1614 ? io_enq_uops_2_exception : rob_exception_2_25));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_26 <=
      ~_GEN_2127
      & (_GEN_69 & _GEN_913 | (_GEN_1615 ? io_enq_uops_2_exception : rob_exception_2_26));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_27 <=
      ~_GEN_2128
      & (_GEN_69 & _GEN_914 | (_GEN_1616 ? io_enq_uops_2_exception : rob_exception_2_27));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_28 <=
      ~_GEN_2129
      & (_GEN_69 & _GEN_915 | (_GEN_1617 ? io_enq_uops_2_exception : rob_exception_2_28));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_29 <=
      ~_GEN_2130
      & (_GEN_69 & _GEN_916 | (_GEN_1618 ? io_enq_uops_2_exception : rob_exception_2_29));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_30 <=
      ~_GEN_2131
      & (_GEN_69 & _GEN_917 | (_GEN_1619 ? io_enq_uops_2_exception : rob_exception_2_30));	// rob.scala:307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_exception_2_31 <=
      ~_GEN_2132
      & (_GEN_69 & (&(io_lxcpt_bits_uop_rob_idx[6:2]))
         | (_GEN_1620 ? io_enq_uops_2_exception : rob_exception_2_31));	// rob.scala:236:31, :268:25, :307:32, :311:28, :323:29, :324:31, :329:31, :390:{26,79}, :391:59, :433:20, :434:30, :435:30
    rob_predicated_2_0 <=
      ~(_GEN_65 & _GEN_666)
      & (_GEN_1941
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_476 | _GEN_1813 | _GEN_61 & _GEN_286)
             & (_GEN_1685
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1589 & rob_predicated_2_0));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_1 <=
      ~(_GEN_65 & _GEN_669)
      & (_GEN_1942
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_479 | _GEN_1814 | _GEN_61 & _GEN_289)
             & (_GEN_1686
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1590 & rob_predicated_2_1));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_2 <=
      ~(_GEN_65 & _GEN_672)
      & (_GEN_1943
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_482 | _GEN_1815 | _GEN_61 & _GEN_292)
             & (_GEN_1687
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1591 & rob_predicated_2_2));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_3 <=
      ~(_GEN_65 & _GEN_675)
      & (_GEN_1944
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_485 | _GEN_1816 | _GEN_61 & _GEN_295)
             & (_GEN_1688
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1592 & rob_predicated_2_3));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_4 <=
      ~(_GEN_65 & _GEN_678)
      & (_GEN_1945
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_488 | _GEN_1817 | _GEN_61 & _GEN_298)
             & (_GEN_1689
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1593 & rob_predicated_2_4));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_5 <=
      ~(_GEN_65 & _GEN_681)
      & (_GEN_1946
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_491 | _GEN_1818 | _GEN_61 & _GEN_301)
             & (_GEN_1690
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1594 & rob_predicated_2_5));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_6 <=
      ~(_GEN_65 & _GEN_684)
      & (_GEN_1947
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_494 | _GEN_1819 | _GEN_61 & _GEN_304)
             & (_GEN_1691
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1595 & rob_predicated_2_6));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_7 <=
      ~(_GEN_65 & _GEN_687)
      & (_GEN_1948
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_497 | _GEN_1820 | _GEN_61 & _GEN_307)
             & (_GEN_1692
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1596 & rob_predicated_2_7));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_8 <=
      ~(_GEN_65 & _GEN_690)
      & (_GEN_1949
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_500 | _GEN_1821 | _GEN_61 & _GEN_310)
             & (_GEN_1693
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1597 & rob_predicated_2_8));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_9 <=
      ~(_GEN_65 & _GEN_693)
      & (_GEN_1950
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_503 | _GEN_1822 | _GEN_61 & _GEN_313)
             & (_GEN_1694
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1598 & rob_predicated_2_9));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_10 <=
      ~(_GEN_65 & _GEN_696)
      & (_GEN_1951
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_506 | _GEN_1823 | _GEN_61 & _GEN_316)
             & (_GEN_1695
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1599 & rob_predicated_2_10));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_11 <=
      ~(_GEN_65 & _GEN_699)
      & (_GEN_1952
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_509 | _GEN_1824 | _GEN_61 & _GEN_319)
             & (_GEN_1696
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1600 & rob_predicated_2_11));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_12 <=
      ~(_GEN_65 & _GEN_702)
      & (_GEN_1953
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_512 | _GEN_1825 | _GEN_61 & _GEN_322)
             & (_GEN_1697
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1601 & rob_predicated_2_12));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_13 <=
      ~(_GEN_65 & _GEN_705)
      & (_GEN_1954
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_515 | _GEN_1826 | _GEN_61 & _GEN_325)
             & (_GEN_1698
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1602 & rob_predicated_2_13));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_14 <=
      ~(_GEN_65 & _GEN_708)
      & (_GEN_1955
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_518 | _GEN_1827 | _GEN_61 & _GEN_328)
             & (_GEN_1699
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1603 & rob_predicated_2_14));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_15 <=
      ~(_GEN_65 & _GEN_711)
      & (_GEN_1956
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_521 | _GEN_1828 | _GEN_61 & _GEN_331)
             & (_GEN_1700
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1604 & rob_predicated_2_15));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_16 <=
      ~(_GEN_65 & _GEN_714)
      & (_GEN_1957
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_524 | _GEN_1829 | _GEN_61 & _GEN_334)
             & (_GEN_1701
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1605 & rob_predicated_2_16));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_17 <=
      ~(_GEN_65 & _GEN_717)
      & (_GEN_1958
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_527 | _GEN_1830 | _GEN_61 & _GEN_337)
             & (_GEN_1702
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1606 & rob_predicated_2_17));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_18 <=
      ~(_GEN_65 & _GEN_720)
      & (_GEN_1959
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_530 | _GEN_1831 | _GEN_61 & _GEN_340)
             & (_GEN_1703
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1607 & rob_predicated_2_18));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_19 <=
      ~(_GEN_65 & _GEN_723)
      & (_GEN_1960
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_533 | _GEN_1832 | _GEN_61 & _GEN_343)
             & (_GEN_1704
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1608 & rob_predicated_2_19));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_20 <=
      ~(_GEN_65 & _GEN_726)
      & (_GEN_1961
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_536 | _GEN_1833 | _GEN_61 & _GEN_346)
             & (_GEN_1705
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1609 & rob_predicated_2_20));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_21 <=
      ~(_GEN_65 & _GEN_729)
      & (_GEN_1962
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_539 | _GEN_1834 | _GEN_61 & _GEN_349)
             & (_GEN_1706
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1610 & rob_predicated_2_21));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_22 <=
      ~(_GEN_65 & _GEN_732)
      & (_GEN_1963
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_542 | _GEN_1835 | _GEN_61 & _GEN_352)
             & (_GEN_1707
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1611 & rob_predicated_2_22));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_23 <=
      ~(_GEN_65 & _GEN_735)
      & (_GEN_1964
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_545 | _GEN_1836 | _GEN_61 & _GEN_355)
             & (_GEN_1708
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1612 & rob_predicated_2_23));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_24 <=
      ~(_GEN_65 & _GEN_738)
      & (_GEN_1965
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_548 | _GEN_1837 | _GEN_61 & _GEN_358)
             & (_GEN_1709
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1613 & rob_predicated_2_24));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_25 <=
      ~(_GEN_65 & _GEN_741)
      & (_GEN_1966
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_551 | _GEN_1838 | _GEN_61 & _GEN_361)
             & (_GEN_1710
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1614 & rob_predicated_2_25));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_26 <=
      ~(_GEN_65 & _GEN_744)
      & (_GEN_1967
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_554 | _GEN_1839 | _GEN_61 & _GEN_364)
             & (_GEN_1711
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1615 & rob_predicated_2_26));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_27 <=
      ~(_GEN_65 & _GEN_747)
      & (_GEN_1968
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_557 | _GEN_1840 | _GEN_61 & _GEN_367)
             & (_GEN_1712
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1616 & rob_predicated_2_27));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_28 <=
      ~(_GEN_65 & _GEN_750)
      & (_GEN_1969
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_560 | _GEN_1841 | _GEN_61 & _GEN_370)
             & (_GEN_1713
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1617 & rob_predicated_2_28));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_29 <=
      ~(_GEN_65 & _GEN_753)
      & (_GEN_1970
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_563 | _GEN_1842 | _GEN_61 & _GEN_373)
             & (_GEN_1714
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1618 & rob_predicated_2_29));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_30 <=
      ~(_GEN_65 & _GEN_756)
      & (_GEN_1971
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & _GEN_566 | _GEN_1843 | _GEN_61 & _GEN_376)
             & (_GEN_1715
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1619 & rob_predicated_2_30));	// rob.scala:307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    rob_predicated_2_31 <=
      ~(_GEN_65 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])))
      & (_GEN_1972
           ? io_wb_resps_4_bits_predicated
           : ~(_GEN_63 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1844 | _GEN_61
               & (&(io_wb_resps_1_bits_uop_rob_idx[6:2])))
             & (_GEN_1716
                  ? io_wb_resps_0_bits_predicated
                  : ~_GEN_1620 & rob_predicated_2_31));	// rob.scala:236:31, :268:25, :307:32, :312:29, :323:29, :324:31, :330:34, :346:{27,69}, :347:31, :349:34
    block_commit_REG <= exception_thrown;	// rob.scala:540:94, :545:85
    block_commit_REG_1 <= exception_thrown;	// rob.scala:540:131, :545:85
    block_commit_REG_2 <= block_commit_REG_1;	// rob.scala:540:{123,131}
    REG <= exception_thrown;	// rob.scala:545:85, :808:30
    REG_1 <= REG;	// rob.scala:808:{22,30}
    REG_2 <= exception_thrown;	// rob.scala:545:85, :824:22
    _GEN_2169 =
      {{rob_head_uses_ldq_0},
       {_GEN_81[rob_head]},
       {_GEN_51[rob_head]},
       {rob_head_uses_ldq_0}};	// rob.scala:224:29, :411:25, :484:26, :865:98
    io_com_load_is_at_rob_head_REG <=
      _GEN_2169[rob_head_vals_0 ? 2'h0 : rob_head_vals_1 ? 2'h1 : 2'h2]
      & ~(will_commit_0 | will_commit_1 | will_commit_2);	// Mux.scala:47:69, rob.scala:221:26, :236:31, :398:49, :540:33, :547:70, :865:{40,98}, :866:{41,62}
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:1260];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [10:0] i = 11'h0; i < 11'h4ED; i += 11'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        rob_state = _RANDOM[11'h0][1:0];	// rob.scala:221:26
        rob_head = _RANDOM[11'h0][6:2];	// rob.scala:221:26, :224:29
        rob_head_lsb = _RANDOM[11'h0][8:7];	// rob.scala:221:26, :225:29
        rob_tail = _RANDOM[11'h0][13:9];	// rob.scala:221:26, :228:29
        rob_tail_lsb = _RANDOM[11'h0][15:14];	// rob.scala:221:26, :229:29
        rob_pnr = _RANDOM[11'h0][20:16];	// rob.scala:221:26, :232:29
        rob_pnr_lsb = _RANDOM[11'h0][22:21];	// rob.scala:221:26, :233:29
        maybe_full = _RANDOM[11'h0][23];	// rob.scala:221:26, :239:29
        r_xcpt_val = _RANDOM[11'h0][24];	// rob.scala:221:26, :258:33
        r_xcpt_uop_br_mask = {_RANDOM[11'h5][31:21], _RANDOM[11'h6][4:0]};	// rob.scala:259:29
        r_xcpt_uop_rob_idx = _RANDOM[11'h7][28:22];	// rob.scala:259:29
        r_xcpt_uop_exc_cause =
          {_RANDOM[11'h9][31:22], _RANDOM[11'hA], _RANDOM[11'hB][21:0]};	// rob.scala:259:29
        r_xcpt_badvaddr = {_RANDOM[11'hD][31:19], _RANDOM[11'hE][26:0]};	// rob.scala:260:29
        rob_val_0 = _RANDOM[11'hE][27];	// rob.scala:260:29, :307:32
        rob_val_1 = _RANDOM[11'hE][28];	// rob.scala:260:29, :307:32
        rob_val_2 = _RANDOM[11'hE][29];	// rob.scala:260:29, :307:32
        rob_val_3 = _RANDOM[11'hE][30];	// rob.scala:260:29, :307:32
        rob_val_4 = _RANDOM[11'hE][31];	// rob.scala:260:29, :307:32
        rob_val_5 = _RANDOM[11'hF][0];	// rob.scala:307:32
        rob_val_6 = _RANDOM[11'hF][1];	// rob.scala:307:32
        rob_val_7 = _RANDOM[11'hF][2];	// rob.scala:307:32
        rob_val_8 = _RANDOM[11'hF][3];	// rob.scala:307:32
        rob_val_9 = _RANDOM[11'hF][4];	// rob.scala:307:32
        rob_val_10 = _RANDOM[11'hF][5];	// rob.scala:307:32
        rob_val_11 = _RANDOM[11'hF][6];	// rob.scala:307:32
        rob_val_12 = _RANDOM[11'hF][7];	// rob.scala:307:32
        rob_val_13 = _RANDOM[11'hF][8];	// rob.scala:307:32
        rob_val_14 = _RANDOM[11'hF][9];	// rob.scala:307:32
        rob_val_15 = _RANDOM[11'hF][10];	// rob.scala:307:32
        rob_val_16 = _RANDOM[11'hF][11];	// rob.scala:307:32
        rob_val_17 = _RANDOM[11'hF][12];	// rob.scala:307:32
        rob_val_18 = _RANDOM[11'hF][13];	// rob.scala:307:32
        rob_val_19 = _RANDOM[11'hF][14];	// rob.scala:307:32
        rob_val_20 = _RANDOM[11'hF][15];	// rob.scala:307:32
        rob_val_21 = _RANDOM[11'hF][16];	// rob.scala:307:32
        rob_val_22 = _RANDOM[11'hF][17];	// rob.scala:307:32
        rob_val_23 = _RANDOM[11'hF][18];	// rob.scala:307:32
        rob_val_24 = _RANDOM[11'hF][19];	// rob.scala:307:32
        rob_val_25 = _RANDOM[11'hF][20];	// rob.scala:307:32
        rob_val_26 = _RANDOM[11'hF][21];	// rob.scala:307:32
        rob_val_27 = _RANDOM[11'hF][22];	// rob.scala:307:32
        rob_val_28 = _RANDOM[11'hF][23];	// rob.scala:307:32
        rob_val_29 = _RANDOM[11'hF][24];	// rob.scala:307:32
        rob_val_30 = _RANDOM[11'hF][25];	// rob.scala:307:32
        rob_val_31 = _RANDOM[11'hF][26];	// rob.scala:307:32
        rob_bsy_0 = _RANDOM[11'hF][27];	// rob.scala:307:32, :308:28
        rob_bsy_1 = _RANDOM[11'hF][28];	// rob.scala:307:32, :308:28
        rob_bsy_2 = _RANDOM[11'hF][29];	// rob.scala:307:32, :308:28
        rob_bsy_3 = _RANDOM[11'hF][30];	// rob.scala:307:32, :308:28
        rob_bsy_4 = _RANDOM[11'hF][31];	// rob.scala:307:32, :308:28
        rob_bsy_5 = _RANDOM[11'h10][0];	// rob.scala:308:28
        rob_bsy_6 = _RANDOM[11'h10][1];	// rob.scala:308:28
        rob_bsy_7 = _RANDOM[11'h10][2];	// rob.scala:308:28
        rob_bsy_8 = _RANDOM[11'h10][3];	// rob.scala:308:28
        rob_bsy_9 = _RANDOM[11'h10][4];	// rob.scala:308:28
        rob_bsy_10 = _RANDOM[11'h10][5];	// rob.scala:308:28
        rob_bsy_11 = _RANDOM[11'h10][6];	// rob.scala:308:28
        rob_bsy_12 = _RANDOM[11'h10][7];	// rob.scala:308:28
        rob_bsy_13 = _RANDOM[11'h10][8];	// rob.scala:308:28
        rob_bsy_14 = _RANDOM[11'h10][9];	// rob.scala:308:28
        rob_bsy_15 = _RANDOM[11'h10][10];	// rob.scala:308:28
        rob_bsy_16 = _RANDOM[11'h10][11];	// rob.scala:308:28
        rob_bsy_17 = _RANDOM[11'h10][12];	// rob.scala:308:28
        rob_bsy_18 = _RANDOM[11'h10][13];	// rob.scala:308:28
        rob_bsy_19 = _RANDOM[11'h10][14];	// rob.scala:308:28
        rob_bsy_20 = _RANDOM[11'h10][15];	// rob.scala:308:28
        rob_bsy_21 = _RANDOM[11'h10][16];	// rob.scala:308:28
        rob_bsy_22 = _RANDOM[11'h10][17];	// rob.scala:308:28
        rob_bsy_23 = _RANDOM[11'h10][18];	// rob.scala:308:28
        rob_bsy_24 = _RANDOM[11'h10][19];	// rob.scala:308:28
        rob_bsy_25 = _RANDOM[11'h10][20];	// rob.scala:308:28
        rob_bsy_26 = _RANDOM[11'h10][21];	// rob.scala:308:28
        rob_bsy_27 = _RANDOM[11'h10][22];	// rob.scala:308:28
        rob_bsy_28 = _RANDOM[11'h10][23];	// rob.scala:308:28
        rob_bsy_29 = _RANDOM[11'h10][24];	// rob.scala:308:28
        rob_bsy_30 = _RANDOM[11'h10][25];	// rob.scala:308:28
        rob_bsy_31 = _RANDOM[11'h10][26];	// rob.scala:308:28
        rob_unsafe_0 = _RANDOM[11'h10][27];	// rob.scala:308:28, :309:28
        rob_unsafe_1 = _RANDOM[11'h10][28];	// rob.scala:308:28, :309:28
        rob_unsafe_2 = _RANDOM[11'h10][29];	// rob.scala:308:28, :309:28
        rob_unsafe_3 = _RANDOM[11'h10][30];	// rob.scala:308:28, :309:28
        rob_unsafe_4 = _RANDOM[11'h10][31];	// rob.scala:308:28, :309:28
        rob_unsafe_5 = _RANDOM[11'h11][0];	// rob.scala:309:28
        rob_unsafe_6 = _RANDOM[11'h11][1];	// rob.scala:309:28
        rob_unsafe_7 = _RANDOM[11'h11][2];	// rob.scala:309:28
        rob_unsafe_8 = _RANDOM[11'h11][3];	// rob.scala:309:28
        rob_unsafe_9 = _RANDOM[11'h11][4];	// rob.scala:309:28
        rob_unsafe_10 = _RANDOM[11'h11][5];	// rob.scala:309:28
        rob_unsafe_11 = _RANDOM[11'h11][6];	// rob.scala:309:28
        rob_unsafe_12 = _RANDOM[11'h11][7];	// rob.scala:309:28
        rob_unsafe_13 = _RANDOM[11'h11][8];	// rob.scala:309:28
        rob_unsafe_14 = _RANDOM[11'h11][9];	// rob.scala:309:28
        rob_unsafe_15 = _RANDOM[11'h11][10];	// rob.scala:309:28
        rob_unsafe_16 = _RANDOM[11'h11][11];	// rob.scala:309:28
        rob_unsafe_17 = _RANDOM[11'h11][12];	// rob.scala:309:28
        rob_unsafe_18 = _RANDOM[11'h11][13];	// rob.scala:309:28
        rob_unsafe_19 = _RANDOM[11'h11][14];	// rob.scala:309:28
        rob_unsafe_20 = _RANDOM[11'h11][15];	// rob.scala:309:28
        rob_unsafe_21 = _RANDOM[11'h11][16];	// rob.scala:309:28
        rob_unsafe_22 = _RANDOM[11'h11][17];	// rob.scala:309:28
        rob_unsafe_23 = _RANDOM[11'h11][18];	// rob.scala:309:28
        rob_unsafe_24 = _RANDOM[11'h11][19];	// rob.scala:309:28
        rob_unsafe_25 = _RANDOM[11'h11][20];	// rob.scala:309:28
        rob_unsafe_26 = _RANDOM[11'h11][21];	// rob.scala:309:28
        rob_unsafe_27 = _RANDOM[11'h11][22];	// rob.scala:309:28
        rob_unsafe_28 = _RANDOM[11'h11][23];	// rob.scala:309:28
        rob_unsafe_29 = _RANDOM[11'h11][24];	// rob.scala:309:28
        rob_unsafe_30 = _RANDOM[11'h11][25];	// rob.scala:309:28
        rob_unsafe_31 = _RANDOM[11'h11][26];	// rob.scala:309:28
        rob_uop_0_uopc = {_RANDOM[11'h11][31:27], _RANDOM[11'h12][1:0]};	// rob.scala:309:28, :310:28
        rob_uop_0_is_rvc = _RANDOM[11'h14][2];	// rob.scala:310:28
        rob_uop_0_br_mask = {_RANDOM[11'h16][31:23], _RANDOM[11'h17][6:0]};	// rob.scala:310:28
        rob_uop_0_ftq_idx = _RANDOM[11'h17][15:11];	// rob.scala:310:28
        rob_uop_0_edge_inst = _RANDOM[11'h17][16];	// rob.scala:310:28
        rob_uop_0_pc_lob = _RANDOM[11'h17][22:17];	// rob.scala:310:28
        rob_uop_0_pdst = _RANDOM[11'h19][17:11];	// rob.scala:310:28
        rob_uop_0_stale_pdst = _RANDOM[11'h1A][22:16];	// rob.scala:310:28
        rob_uop_0_is_fencei = _RANDOM[11'h1D][2];	// rob.scala:310:28
        rob_uop_0_uses_ldq = _RANDOM[11'h1D][4];	// rob.scala:310:28
        rob_uop_0_uses_stq = _RANDOM[11'h1D][5];	// rob.scala:310:28
        rob_uop_0_is_sys_pc2epc = _RANDOM[11'h1D][6];	// rob.scala:310:28
        rob_uop_0_flush_on_commit = _RANDOM[11'h1D][8];	// rob.scala:310:28
        rob_uop_0_ldst = _RANDOM[11'h1D][15:10];	// rob.scala:310:28
        rob_uop_0_ldst_val = _RANDOM[11'h1E][2];	// rob.scala:310:28
        rob_uop_0_dst_rtype = _RANDOM[11'h1E][4:3];	// rob.scala:310:28
        rob_uop_0_fp_val = _RANDOM[11'h1E][10];	// rob.scala:310:28
        rob_uop_1_uopc = _RANDOM[11'h1E][27:21];	// rob.scala:310:28
        rob_uop_1_is_rvc = _RANDOM[11'h20][28];	// rob.scala:310:28
        rob_uop_1_br_mask = {_RANDOM[11'h23][31:17], _RANDOM[11'h24][0]};	// rob.scala:310:28
        rob_uop_1_ftq_idx = _RANDOM[11'h24][9:5];	// rob.scala:310:28
        rob_uop_1_edge_inst = _RANDOM[11'h24][10];	// rob.scala:310:28
        rob_uop_1_pc_lob = _RANDOM[11'h24][16:11];	// rob.scala:310:28
        rob_uop_1_pdst = _RANDOM[11'h26][11:5];	// rob.scala:310:28
        rob_uop_1_stale_pdst = _RANDOM[11'h27][16:10];	// rob.scala:310:28
        rob_uop_1_is_fencei = _RANDOM[11'h29][28];	// rob.scala:310:28
        rob_uop_1_uses_ldq = _RANDOM[11'h29][30];	// rob.scala:310:28
        rob_uop_1_uses_stq = _RANDOM[11'h29][31];	// rob.scala:310:28
        rob_uop_1_is_sys_pc2epc = _RANDOM[11'h2A][0];	// rob.scala:310:28
        rob_uop_1_flush_on_commit = _RANDOM[11'h2A][2];	// rob.scala:310:28
        rob_uop_1_ldst = _RANDOM[11'h2A][9:4];	// rob.scala:310:28
        rob_uop_1_ldst_val = _RANDOM[11'h2A][28];	// rob.scala:310:28
        rob_uop_1_dst_rtype = _RANDOM[11'h2A][30:29];	// rob.scala:310:28
        rob_uop_1_fp_val = _RANDOM[11'h2B][4];	// rob.scala:310:28
        rob_uop_2_uopc = _RANDOM[11'h2B][21:15];	// rob.scala:310:28
        rob_uop_2_is_rvc = _RANDOM[11'h2D][22];	// rob.scala:310:28
        rob_uop_2_br_mask = _RANDOM[11'h30][26:11];	// rob.scala:310:28
        rob_uop_2_ftq_idx = {_RANDOM[11'h30][31], _RANDOM[11'h31][3:0]};	// rob.scala:310:28
        rob_uop_2_edge_inst = _RANDOM[11'h31][4];	// rob.scala:310:28
        rob_uop_2_pc_lob = _RANDOM[11'h31][10:5];	// rob.scala:310:28
        rob_uop_2_pdst = {_RANDOM[11'h32][31], _RANDOM[11'h33][5:0]};	// rob.scala:310:28
        rob_uop_2_stale_pdst = _RANDOM[11'h34][10:4];	// rob.scala:310:28
        rob_uop_2_is_fencei = _RANDOM[11'h36][22];	// rob.scala:310:28
        rob_uop_2_uses_ldq = _RANDOM[11'h36][24];	// rob.scala:310:28
        rob_uop_2_uses_stq = _RANDOM[11'h36][25];	// rob.scala:310:28
        rob_uop_2_is_sys_pc2epc = _RANDOM[11'h36][26];	// rob.scala:310:28
        rob_uop_2_flush_on_commit = _RANDOM[11'h36][28];	// rob.scala:310:28
        rob_uop_2_ldst = {_RANDOM[11'h36][31:30], _RANDOM[11'h37][3:0]};	// rob.scala:310:28
        rob_uop_2_ldst_val = _RANDOM[11'h37][22];	// rob.scala:310:28
        rob_uop_2_dst_rtype = _RANDOM[11'h37][24:23];	// rob.scala:310:28
        rob_uop_2_fp_val = _RANDOM[11'h37][30];	// rob.scala:310:28
        rob_uop_3_uopc = _RANDOM[11'h38][15:9];	// rob.scala:310:28
        rob_uop_3_is_rvc = _RANDOM[11'h3A][16];	// rob.scala:310:28
        rob_uop_3_br_mask = _RANDOM[11'h3D][20:5];	// rob.scala:310:28
        rob_uop_3_ftq_idx = _RANDOM[11'h3D][29:25];	// rob.scala:310:28
        rob_uop_3_edge_inst = _RANDOM[11'h3D][30];	// rob.scala:310:28
        rob_uop_3_pc_lob = {_RANDOM[11'h3D][31], _RANDOM[11'h3E][4:0]};	// rob.scala:310:28
        rob_uop_3_pdst = _RANDOM[11'h3F][31:25];	// rob.scala:310:28
        rob_uop_3_stale_pdst = {_RANDOM[11'h40][31:30], _RANDOM[11'h41][4:0]};	// rob.scala:310:28
        rob_uop_3_is_fencei = _RANDOM[11'h43][16];	// rob.scala:310:28
        rob_uop_3_uses_ldq = _RANDOM[11'h43][18];	// rob.scala:310:28
        rob_uop_3_uses_stq = _RANDOM[11'h43][19];	// rob.scala:310:28
        rob_uop_3_is_sys_pc2epc = _RANDOM[11'h43][20];	// rob.scala:310:28
        rob_uop_3_flush_on_commit = _RANDOM[11'h43][22];	// rob.scala:310:28
        rob_uop_3_ldst = _RANDOM[11'h43][29:24];	// rob.scala:310:28
        rob_uop_3_ldst_val = _RANDOM[11'h44][16];	// rob.scala:310:28
        rob_uop_3_dst_rtype = _RANDOM[11'h44][18:17];	// rob.scala:310:28
        rob_uop_3_fp_val = _RANDOM[11'h44][24];	// rob.scala:310:28
        rob_uop_4_uopc = _RANDOM[11'h45][9:3];	// rob.scala:310:28
        rob_uop_4_is_rvc = _RANDOM[11'h47][10];	// rob.scala:310:28
        rob_uop_4_br_mask = {_RANDOM[11'h49][31], _RANDOM[11'h4A][14:0]};	// rob.scala:310:28
        rob_uop_4_ftq_idx = _RANDOM[11'h4A][23:19];	// rob.scala:310:28
        rob_uop_4_edge_inst = _RANDOM[11'h4A][24];	// rob.scala:310:28
        rob_uop_4_pc_lob = _RANDOM[11'h4A][30:25];	// rob.scala:310:28
        rob_uop_4_pdst = _RANDOM[11'h4C][25:19];	// rob.scala:310:28
        rob_uop_4_stale_pdst = _RANDOM[11'h4D][30:24];	// rob.scala:310:28
        rob_uop_4_is_fencei = _RANDOM[11'h50][10];	// rob.scala:310:28
        rob_uop_4_uses_ldq = _RANDOM[11'h50][12];	// rob.scala:310:28
        rob_uop_4_uses_stq = _RANDOM[11'h50][13];	// rob.scala:310:28
        rob_uop_4_is_sys_pc2epc = _RANDOM[11'h50][14];	// rob.scala:310:28
        rob_uop_4_flush_on_commit = _RANDOM[11'h50][16];	// rob.scala:310:28
        rob_uop_4_ldst = _RANDOM[11'h50][23:18];	// rob.scala:310:28
        rob_uop_4_ldst_val = _RANDOM[11'h51][10];	// rob.scala:310:28
        rob_uop_4_dst_rtype = _RANDOM[11'h51][12:11];	// rob.scala:310:28
        rob_uop_4_fp_val = _RANDOM[11'h51][18];	// rob.scala:310:28
        rob_uop_5_uopc = {_RANDOM[11'h51][31:29], _RANDOM[11'h52][3:0]};	// rob.scala:310:28
        rob_uop_5_is_rvc = _RANDOM[11'h54][4];	// rob.scala:310:28
        rob_uop_5_br_mask = {_RANDOM[11'h56][31:25], _RANDOM[11'h57][8:0]};	// rob.scala:310:28
        rob_uop_5_ftq_idx = _RANDOM[11'h57][17:13];	// rob.scala:310:28
        rob_uop_5_edge_inst = _RANDOM[11'h57][18];	// rob.scala:310:28
        rob_uop_5_pc_lob = _RANDOM[11'h57][24:19];	// rob.scala:310:28
        rob_uop_5_pdst = _RANDOM[11'h59][19:13];	// rob.scala:310:28
        rob_uop_5_stale_pdst = _RANDOM[11'h5A][24:18];	// rob.scala:310:28
        rob_uop_5_is_fencei = _RANDOM[11'h5D][4];	// rob.scala:310:28
        rob_uop_5_uses_ldq = _RANDOM[11'h5D][6];	// rob.scala:310:28
        rob_uop_5_uses_stq = _RANDOM[11'h5D][7];	// rob.scala:310:28
        rob_uop_5_is_sys_pc2epc = _RANDOM[11'h5D][8];	// rob.scala:310:28
        rob_uop_5_flush_on_commit = _RANDOM[11'h5D][10];	// rob.scala:310:28
        rob_uop_5_ldst = _RANDOM[11'h5D][17:12];	// rob.scala:310:28
        rob_uop_5_ldst_val = _RANDOM[11'h5E][4];	// rob.scala:310:28
        rob_uop_5_dst_rtype = _RANDOM[11'h5E][6:5];	// rob.scala:310:28
        rob_uop_5_fp_val = _RANDOM[11'h5E][12];	// rob.scala:310:28
        rob_uop_6_uopc = _RANDOM[11'h5E][29:23];	// rob.scala:310:28
        rob_uop_6_is_rvc = _RANDOM[11'h60][30];	// rob.scala:310:28
        rob_uop_6_br_mask = {_RANDOM[11'h63][31:19], _RANDOM[11'h64][2:0]};	// rob.scala:310:28
        rob_uop_6_ftq_idx = _RANDOM[11'h64][11:7];	// rob.scala:310:28
        rob_uop_6_edge_inst = _RANDOM[11'h64][12];	// rob.scala:310:28
        rob_uop_6_pc_lob = _RANDOM[11'h64][18:13];	// rob.scala:310:28
        rob_uop_6_pdst = _RANDOM[11'h66][13:7];	// rob.scala:310:28
        rob_uop_6_stale_pdst = _RANDOM[11'h67][18:12];	// rob.scala:310:28
        rob_uop_6_is_fencei = _RANDOM[11'h69][30];	// rob.scala:310:28
        rob_uop_6_uses_ldq = _RANDOM[11'h6A][0];	// rob.scala:310:28
        rob_uop_6_uses_stq = _RANDOM[11'h6A][1];	// rob.scala:310:28
        rob_uop_6_is_sys_pc2epc = _RANDOM[11'h6A][2];	// rob.scala:310:28
        rob_uop_6_flush_on_commit = _RANDOM[11'h6A][4];	// rob.scala:310:28
        rob_uop_6_ldst = _RANDOM[11'h6A][11:6];	// rob.scala:310:28
        rob_uop_6_ldst_val = _RANDOM[11'h6A][30];	// rob.scala:310:28
        rob_uop_6_dst_rtype = {_RANDOM[11'h6A][31], _RANDOM[11'h6B][0]};	// rob.scala:310:28
        rob_uop_6_fp_val = _RANDOM[11'h6B][6];	// rob.scala:310:28
        rob_uop_7_uopc = _RANDOM[11'h6B][23:17];	// rob.scala:310:28
        rob_uop_7_is_rvc = _RANDOM[11'h6D][24];	// rob.scala:310:28
        rob_uop_7_br_mask = _RANDOM[11'h70][28:13];	// rob.scala:310:28
        rob_uop_7_ftq_idx = _RANDOM[11'h71][5:1];	// rob.scala:310:28
        rob_uop_7_edge_inst = _RANDOM[11'h71][6];	// rob.scala:310:28
        rob_uop_7_pc_lob = _RANDOM[11'h71][12:7];	// rob.scala:310:28
        rob_uop_7_pdst = _RANDOM[11'h73][7:1];	// rob.scala:310:28
        rob_uop_7_stale_pdst = _RANDOM[11'h74][12:6];	// rob.scala:310:28
        rob_uop_7_is_fencei = _RANDOM[11'h76][24];	// rob.scala:310:28
        rob_uop_7_uses_ldq = _RANDOM[11'h76][26];	// rob.scala:310:28
        rob_uop_7_uses_stq = _RANDOM[11'h76][27];	// rob.scala:310:28
        rob_uop_7_is_sys_pc2epc = _RANDOM[11'h76][28];	// rob.scala:310:28
        rob_uop_7_flush_on_commit = _RANDOM[11'h76][30];	// rob.scala:310:28
        rob_uop_7_ldst = _RANDOM[11'h77][5:0];	// rob.scala:310:28
        rob_uop_7_ldst_val = _RANDOM[11'h77][24];	// rob.scala:310:28
        rob_uop_7_dst_rtype = _RANDOM[11'h77][26:25];	// rob.scala:310:28
        rob_uop_7_fp_val = _RANDOM[11'h78][0];	// rob.scala:310:28
        rob_uop_8_uopc = _RANDOM[11'h78][17:11];	// rob.scala:310:28
        rob_uop_8_is_rvc = _RANDOM[11'h7A][18];	// rob.scala:310:28
        rob_uop_8_br_mask = _RANDOM[11'h7D][22:7];	// rob.scala:310:28
        rob_uop_8_ftq_idx = _RANDOM[11'h7D][31:27];	// rob.scala:310:28
        rob_uop_8_edge_inst = _RANDOM[11'h7E][0];	// rob.scala:310:28
        rob_uop_8_pc_lob = _RANDOM[11'h7E][6:1];	// rob.scala:310:28
        rob_uop_8_pdst = {_RANDOM[11'h7F][31:27], _RANDOM[11'h80][1:0]};	// rob.scala:310:28
        rob_uop_8_stale_pdst = _RANDOM[11'h81][6:0];	// rob.scala:310:28
        rob_uop_8_is_fencei = _RANDOM[11'h83][18];	// rob.scala:310:28
        rob_uop_8_uses_ldq = _RANDOM[11'h83][20];	// rob.scala:310:28
        rob_uop_8_uses_stq = _RANDOM[11'h83][21];	// rob.scala:310:28
        rob_uop_8_is_sys_pc2epc = _RANDOM[11'h83][22];	// rob.scala:310:28
        rob_uop_8_flush_on_commit = _RANDOM[11'h83][24];	// rob.scala:310:28
        rob_uop_8_ldst = _RANDOM[11'h83][31:26];	// rob.scala:310:28
        rob_uop_8_ldst_val = _RANDOM[11'h84][18];	// rob.scala:310:28
        rob_uop_8_dst_rtype = _RANDOM[11'h84][20:19];	// rob.scala:310:28
        rob_uop_8_fp_val = _RANDOM[11'h84][26];	// rob.scala:310:28
        rob_uop_9_uopc = _RANDOM[11'h85][11:5];	// rob.scala:310:28
        rob_uop_9_is_rvc = _RANDOM[11'h87][12];	// rob.scala:310:28
        rob_uop_9_br_mask = _RANDOM[11'h8A][16:1];	// rob.scala:310:28
        rob_uop_9_ftq_idx = _RANDOM[11'h8A][25:21];	// rob.scala:310:28
        rob_uop_9_edge_inst = _RANDOM[11'h8A][26];	// rob.scala:310:28
        rob_uop_9_pc_lob = {_RANDOM[11'h8A][31:27], _RANDOM[11'h8B][0]};	// rob.scala:310:28
        rob_uop_9_pdst = _RANDOM[11'h8C][27:21];	// rob.scala:310:28
        rob_uop_9_stale_pdst = {_RANDOM[11'h8D][31:26], _RANDOM[11'h8E][0]};	// rob.scala:310:28
        rob_uop_9_is_fencei = _RANDOM[11'h90][12];	// rob.scala:310:28
        rob_uop_9_uses_ldq = _RANDOM[11'h90][14];	// rob.scala:310:28
        rob_uop_9_uses_stq = _RANDOM[11'h90][15];	// rob.scala:310:28
        rob_uop_9_is_sys_pc2epc = _RANDOM[11'h90][16];	// rob.scala:310:28
        rob_uop_9_flush_on_commit = _RANDOM[11'h90][18];	// rob.scala:310:28
        rob_uop_9_ldst = _RANDOM[11'h90][25:20];	// rob.scala:310:28
        rob_uop_9_ldst_val = _RANDOM[11'h91][12];	// rob.scala:310:28
        rob_uop_9_dst_rtype = _RANDOM[11'h91][14:13];	// rob.scala:310:28
        rob_uop_9_fp_val = _RANDOM[11'h91][20];	// rob.scala:310:28
        rob_uop_10_uopc = {_RANDOM[11'h91][31], _RANDOM[11'h92][5:0]};	// rob.scala:310:28
        rob_uop_10_is_rvc = _RANDOM[11'h94][6];	// rob.scala:310:28
        rob_uop_10_br_mask = {_RANDOM[11'h96][31:27], _RANDOM[11'h97][10:0]};	// rob.scala:310:28
        rob_uop_10_ftq_idx = _RANDOM[11'h97][19:15];	// rob.scala:310:28
        rob_uop_10_edge_inst = _RANDOM[11'h97][20];	// rob.scala:310:28
        rob_uop_10_pc_lob = _RANDOM[11'h97][26:21];	// rob.scala:310:28
        rob_uop_10_pdst = _RANDOM[11'h99][21:15];	// rob.scala:310:28
        rob_uop_10_stale_pdst = _RANDOM[11'h9A][26:20];	// rob.scala:310:28
        rob_uop_10_is_fencei = _RANDOM[11'h9D][6];	// rob.scala:310:28
        rob_uop_10_uses_ldq = _RANDOM[11'h9D][8];	// rob.scala:310:28
        rob_uop_10_uses_stq = _RANDOM[11'h9D][9];	// rob.scala:310:28
        rob_uop_10_is_sys_pc2epc = _RANDOM[11'h9D][10];	// rob.scala:310:28
        rob_uop_10_flush_on_commit = _RANDOM[11'h9D][12];	// rob.scala:310:28
        rob_uop_10_ldst = _RANDOM[11'h9D][19:14];	// rob.scala:310:28
        rob_uop_10_ldst_val = _RANDOM[11'h9E][6];	// rob.scala:310:28
        rob_uop_10_dst_rtype = _RANDOM[11'h9E][8:7];	// rob.scala:310:28
        rob_uop_10_fp_val = _RANDOM[11'h9E][14];	// rob.scala:310:28
        rob_uop_11_uopc = _RANDOM[11'h9E][31:25];	// rob.scala:310:28
        rob_uop_11_is_rvc = _RANDOM[11'hA1][0];	// rob.scala:310:28
        rob_uop_11_br_mask = {_RANDOM[11'hA3][31:21], _RANDOM[11'hA4][4:0]};	// rob.scala:310:28
        rob_uop_11_ftq_idx = _RANDOM[11'hA4][13:9];	// rob.scala:310:28
        rob_uop_11_edge_inst = _RANDOM[11'hA4][14];	// rob.scala:310:28
        rob_uop_11_pc_lob = _RANDOM[11'hA4][20:15];	// rob.scala:310:28
        rob_uop_11_pdst = _RANDOM[11'hA6][15:9];	// rob.scala:310:28
        rob_uop_11_stale_pdst = _RANDOM[11'hA7][20:14];	// rob.scala:310:28
        rob_uop_11_is_fencei = _RANDOM[11'hAA][0];	// rob.scala:310:28
        rob_uop_11_uses_ldq = _RANDOM[11'hAA][2];	// rob.scala:310:28
        rob_uop_11_uses_stq = _RANDOM[11'hAA][3];	// rob.scala:310:28
        rob_uop_11_is_sys_pc2epc = _RANDOM[11'hAA][4];	// rob.scala:310:28
        rob_uop_11_flush_on_commit = _RANDOM[11'hAA][6];	// rob.scala:310:28
        rob_uop_11_ldst = _RANDOM[11'hAA][13:8];	// rob.scala:310:28
        rob_uop_11_ldst_val = _RANDOM[11'hAB][0];	// rob.scala:310:28
        rob_uop_11_dst_rtype = _RANDOM[11'hAB][2:1];	// rob.scala:310:28
        rob_uop_11_fp_val = _RANDOM[11'hAB][8];	// rob.scala:310:28
        rob_uop_12_uopc = _RANDOM[11'hAB][25:19];	// rob.scala:310:28
        rob_uop_12_is_rvc = _RANDOM[11'hAD][26];	// rob.scala:310:28
        rob_uop_12_br_mask = _RANDOM[11'hB0][30:15];	// rob.scala:310:28
        rob_uop_12_ftq_idx = _RANDOM[11'hB1][7:3];	// rob.scala:310:28
        rob_uop_12_edge_inst = _RANDOM[11'hB1][8];	// rob.scala:310:28
        rob_uop_12_pc_lob = _RANDOM[11'hB1][14:9];	// rob.scala:310:28
        rob_uop_12_pdst = _RANDOM[11'hB3][9:3];	// rob.scala:310:28
        rob_uop_12_stale_pdst = _RANDOM[11'hB4][14:8];	// rob.scala:310:28
        rob_uop_12_is_fencei = _RANDOM[11'hB6][26];	// rob.scala:310:28
        rob_uop_12_uses_ldq = _RANDOM[11'hB6][28];	// rob.scala:310:28
        rob_uop_12_uses_stq = _RANDOM[11'hB6][29];	// rob.scala:310:28
        rob_uop_12_is_sys_pc2epc = _RANDOM[11'hB6][30];	// rob.scala:310:28
        rob_uop_12_flush_on_commit = _RANDOM[11'hB7][0];	// rob.scala:310:28
        rob_uop_12_ldst = _RANDOM[11'hB7][7:2];	// rob.scala:310:28
        rob_uop_12_ldst_val = _RANDOM[11'hB7][26];	// rob.scala:310:28
        rob_uop_12_dst_rtype = _RANDOM[11'hB7][28:27];	// rob.scala:310:28
        rob_uop_12_fp_val = _RANDOM[11'hB8][2];	// rob.scala:310:28
        rob_uop_13_uopc = _RANDOM[11'hB8][19:13];	// rob.scala:310:28
        rob_uop_13_is_rvc = _RANDOM[11'hBA][20];	// rob.scala:310:28
        rob_uop_13_br_mask = _RANDOM[11'hBD][24:9];	// rob.scala:310:28
        rob_uop_13_ftq_idx = {_RANDOM[11'hBD][31:29], _RANDOM[11'hBE][1:0]};	// rob.scala:310:28
        rob_uop_13_edge_inst = _RANDOM[11'hBE][2];	// rob.scala:310:28
        rob_uop_13_pc_lob = _RANDOM[11'hBE][8:3];	// rob.scala:310:28
        rob_uop_13_pdst = {_RANDOM[11'hBF][31:29], _RANDOM[11'hC0][3:0]};	// rob.scala:310:28
        rob_uop_13_stale_pdst = _RANDOM[11'hC1][8:2];	// rob.scala:310:28
        rob_uop_13_is_fencei = _RANDOM[11'hC3][20];	// rob.scala:310:28
        rob_uop_13_uses_ldq = _RANDOM[11'hC3][22];	// rob.scala:310:28
        rob_uop_13_uses_stq = _RANDOM[11'hC3][23];	// rob.scala:310:28
        rob_uop_13_is_sys_pc2epc = _RANDOM[11'hC3][24];	// rob.scala:310:28
        rob_uop_13_flush_on_commit = _RANDOM[11'hC3][26];	// rob.scala:310:28
        rob_uop_13_ldst = {_RANDOM[11'hC3][31:28], _RANDOM[11'hC4][1:0]};	// rob.scala:310:28
        rob_uop_13_ldst_val = _RANDOM[11'hC4][20];	// rob.scala:310:28
        rob_uop_13_dst_rtype = _RANDOM[11'hC4][22:21];	// rob.scala:310:28
        rob_uop_13_fp_val = _RANDOM[11'hC4][28];	// rob.scala:310:28
        rob_uop_14_uopc = _RANDOM[11'hC5][13:7];	// rob.scala:310:28
        rob_uop_14_is_rvc = _RANDOM[11'hC7][14];	// rob.scala:310:28
        rob_uop_14_br_mask = _RANDOM[11'hCA][18:3];	// rob.scala:310:28
        rob_uop_14_ftq_idx = _RANDOM[11'hCA][27:23];	// rob.scala:310:28
        rob_uop_14_edge_inst = _RANDOM[11'hCA][28];	// rob.scala:310:28
        rob_uop_14_pc_lob = {_RANDOM[11'hCA][31:29], _RANDOM[11'hCB][2:0]};	// rob.scala:310:28
        rob_uop_14_pdst = _RANDOM[11'hCC][29:23];	// rob.scala:310:28
        rob_uop_14_stale_pdst = {_RANDOM[11'hCD][31:28], _RANDOM[11'hCE][2:0]};	// rob.scala:310:28
        rob_uop_14_is_fencei = _RANDOM[11'hD0][14];	// rob.scala:310:28
        rob_uop_14_uses_ldq = _RANDOM[11'hD0][16];	// rob.scala:310:28
        rob_uop_14_uses_stq = _RANDOM[11'hD0][17];	// rob.scala:310:28
        rob_uop_14_is_sys_pc2epc = _RANDOM[11'hD0][18];	// rob.scala:310:28
        rob_uop_14_flush_on_commit = _RANDOM[11'hD0][20];	// rob.scala:310:28
        rob_uop_14_ldst = _RANDOM[11'hD0][27:22];	// rob.scala:310:28
        rob_uop_14_ldst_val = _RANDOM[11'hD1][14];	// rob.scala:310:28
        rob_uop_14_dst_rtype = _RANDOM[11'hD1][16:15];	// rob.scala:310:28
        rob_uop_14_fp_val = _RANDOM[11'hD1][22];	// rob.scala:310:28
        rob_uop_15_uopc = _RANDOM[11'hD2][7:1];	// rob.scala:310:28
        rob_uop_15_is_rvc = _RANDOM[11'hD4][8];	// rob.scala:310:28
        rob_uop_15_br_mask = {_RANDOM[11'hD6][31:29], _RANDOM[11'hD7][12:0]};	// rob.scala:310:28
        rob_uop_15_ftq_idx = _RANDOM[11'hD7][21:17];	// rob.scala:310:28
        rob_uop_15_edge_inst = _RANDOM[11'hD7][22];	// rob.scala:310:28
        rob_uop_15_pc_lob = _RANDOM[11'hD7][28:23];	// rob.scala:310:28
        rob_uop_15_pdst = _RANDOM[11'hD9][23:17];	// rob.scala:310:28
        rob_uop_15_stale_pdst = _RANDOM[11'hDA][28:22];	// rob.scala:310:28
        rob_uop_15_is_fencei = _RANDOM[11'hDD][8];	// rob.scala:310:28
        rob_uop_15_uses_ldq = _RANDOM[11'hDD][10];	// rob.scala:310:28
        rob_uop_15_uses_stq = _RANDOM[11'hDD][11];	// rob.scala:310:28
        rob_uop_15_is_sys_pc2epc = _RANDOM[11'hDD][12];	// rob.scala:310:28
        rob_uop_15_flush_on_commit = _RANDOM[11'hDD][14];	// rob.scala:310:28
        rob_uop_15_ldst = _RANDOM[11'hDD][21:16];	// rob.scala:310:28
        rob_uop_15_ldst_val = _RANDOM[11'hDE][8];	// rob.scala:310:28
        rob_uop_15_dst_rtype = _RANDOM[11'hDE][10:9];	// rob.scala:310:28
        rob_uop_15_fp_val = _RANDOM[11'hDE][16];	// rob.scala:310:28
        rob_uop_16_uopc = {_RANDOM[11'hDE][31:27], _RANDOM[11'hDF][1:0]};	// rob.scala:310:28
        rob_uop_16_is_rvc = _RANDOM[11'hE1][2];	// rob.scala:310:28
        rob_uop_16_br_mask = {_RANDOM[11'hE3][31:23], _RANDOM[11'hE4][6:0]};	// rob.scala:310:28
        rob_uop_16_ftq_idx = _RANDOM[11'hE4][15:11];	// rob.scala:310:28
        rob_uop_16_edge_inst = _RANDOM[11'hE4][16];	// rob.scala:310:28
        rob_uop_16_pc_lob = _RANDOM[11'hE4][22:17];	// rob.scala:310:28
        rob_uop_16_pdst = _RANDOM[11'hE6][17:11];	// rob.scala:310:28
        rob_uop_16_stale_pdst = _RANDOM[11'hE7][22:16];	// rob.scala:310:28
        rob_uop_16_is_fencei = _RANDOM[11'hEA][2];	// rob.scala:310:28
        rob_uop_16_uses_ldq = _RANDOM[11'hEA][4];	// rob.scala:310:28
        rob_uop_16_uses_stq = _RANDOM[11'hEA][5];	// rob.scala:310:28
        rob_uop_16_is_sys_pc2epc = _RANDOM[11'hEA][6];	// rob.scala:310:28
        rob_uop_16_flush_on_commit = _RANDOM[11'hEA][8];	// rob.scala:310:28
        rob_uop_16_ldst = _RANDOM[11'hEA][15:10];	// rob.scala:310:28
        rob_uop_16_ldst_val = _RANDOM[11'hEB][2];	// rob.scala:310:28
        rob_uop_16_dst_rtype = _RANDOM[11'hEB][4:3];	// rob.scala:310:28
        rob_uop_16_fp_val = _RANDOM[11'hEB][10];	// rob.scala:310:28
        rob_uop_17_uopc = _RANDOM[11'hEB][27:21];	// rob.scala:310:28
        rob_uop_17_is_rvc = _RANDOM[11'hED][28];	// rob.scala:310:28
        rob_uop_17_br_mask = {_RANDOM[11'hF0][31:17], _RANDOM[11'hF1][0]};	// rob.scala:310:28
        rob_uop_17_ftq_idx = _RANDOM[11'hF1][9:5];	// rob.scala:310:28
        rob_uop_17_edge_inst = _RANDOM[11'hF1][10];	// rob.scala:310:28
        rob_uop_17_pc_lob = _RANDOM[11'hF1][16:11];	// rob.scala:310:28
        rob_uop_17_pdst = _RANDOM[11'hF3][11:5];	// rob.scala:310:28
        rob_uop_17_stale_pdst = _RANDOM[11'hF4][16:10];	// rob.scala:310:28
        rob_uop_17_is_fencei = _RANDOM[11'hF6][28];	// rob.scala:310:28
        rob_uop_17_uses_ldq = _RANDOM[11'hF6][30];	// rob.scala:310:28
        rob_uop_17_uses_stq = _RANDOM[11'hF6][31];	// rob.scala:310:28
        rob_uop_17_is_sys_pc2epc = _RANDOM[11'hF7][0];	// rob.scala:310:28
        rob_uop_17_flush_on_commit = _RANDOM[11'hF7][2];	// rob.scala:310:28
        rob_uop_17_ldst = _RANDOM[11'hF7][9:4];	// rob.scala:310:28
        rob_uop_17_ldst_val = _RANDOM[11'hF7][28];	// rob.scala:310:28
        rob_uop_17_dst_rtype = _RANDOM[11'hF7][30:29];	// rob.scala:310:28
        rob_uop_17_fp_val = _RANDOM[11'hF8][4];	// rob.scala:310:28
        rob_uop_18_uopc = _RANDOM[11'hF8][21:15];	// rob.scala:310:28
        rob_uop_18_is_rvc = _RANDOM[11'hFA][22];	// rob.scala:310:28
        rob_uop_18_br_mask = _RANDOM[11'hFD][26:11];	// rob.scala:310:28
        rob_uop_18_ftq_idx = {_RANDOM[11'hFD][31], _RANDOM[11'hFE][3:0]};	// rob.scala:310:28
        rob_uop_18_edge_inst = _RANDOM[11'hFE][4];	// rob.scala:310:28
        rob_uop_18_pc_lob = _RANDOM[11'hFE][10:5];	// rob.scala:310:28
        rob_uop_18_pdst = {_RANDOM[11'hFF][31], _RANDOM[11'h100][5:0]};	// rob.scala:310:28
        rob_uop_18_stale_pdst = _RANDOM[11'h101][10:4];	// rob.scala:310:28
        rob_uop_18_is_fencei = _RANDOM[11'h103][22];	// rob.scala:310:28
        rob_uop_18_uses_ldq = _RANDOM[11'h103][24];	// rob.scala:310:28
        rob_uop_18_uses_stq = _RANDOM[11'h103][25];	// rob.scala:310:28
        rob_uop_18_is_sys_pc2epc = _RANDOM[11'h103][26];	// rob.scala:310:28
        rob_uop_18_flush_on_commit = _RANDOM[11'h103][28];	// rob.scala:310:28
        rob_uop_18_ldst = {_RANDOM[11'h103][31:30], _RANDOM[11'h104][3:0]};	// rob.scala:310:28
        rob_uop_18_ldst_val = _RANDOM[11'h104][22];	// rob.scala:310:28
        rob_uop_18_dst_rtype = _RANDOM[11'h104][24:23];	// rob.scala:310:28
        rob_uop_18_fp_val = _RANDOM[11'h104][30];	// rob.scala:310:28
        rob_uop_19_uopc = _RANDOM[11'h105][15:9];	// rob.scala:310:28
        rob_uop_19_is_rvc = _RANDOM[11'h107][16];	// rob.scala:310:28
        rob_uop_19_br_mask = _RANDOM[11'h10A][20:5];	// rob.scala:310:28
        rob_uop_19_ftq_idx = _RANDOM[11'h10A][29:25];	// rob.scala:310:28
        rob_uop_19_edge_inst = _RANDOM[11'h10A][30];	// rob.scala:310:28
        rob_uop_19_pc_lob = {_RANDOM[11'h10A][31], _RANDOM[11'h10B][4:0]};	// rob.scala:310:28
        rob_uop_19_pdst = _RANDOM[11'h10C][31:25];	// rob.scala:310:28
        rob_uop_19_stale_pdst = {_RANDOM[11'h10D][31:30], _RANDOM[11'h10E][4:0]};	// rob.scala:310:28
        rob_uop_19_is_fencei = _RANDOM[11'h110][16];	// rob.scala:310:28
        rob_uop_19_uses_ldq = _RANDOM[11'h110][18];	// rob.scala:310:28
        rob_uop_19_uses_stq = _RANDOM[11'h110][19];	// rob.scala:310:28
        rob_uop_19_is_sys_pc2epc = _RANDOM[11'h110][20];	// rob.scala:310:28
        rob_uop_19_flush_on_commit = _RANDOM[11'h110][22];	// rob.scala:310:28
        rob_uop_19_ldst = _RANDOM[11'h110][29:24];	// rob.scala:310:28
        rob_uop_19_ldst_val = _RANDOM[11'h111][16];	// rob.scala:310:28
        rob_uop_19_dst_rtype = _RANDOM[11'h111][18:17];	// rob.scala:310:28
        rob_uop_19_fp_val = _RANDOM[11'h111][24];	// rob.scala:310:28
        rob_uop_20_uopc = _RANDOM[11'h112][9:3];	// rob.scala:310:28
        rob_uop_20_is_rvc = _RANDOM[11'h114][10];	// rob.scala:310:28
        rob_uop_20_br_mask = {_RANDOM[11'h116][31], _RANDOM[11'h117][14:0]};	// rob.scala:310:28
        rob_uop_20_ftq_idx = _RANDOM[11'h117][23:19];	// rob.scala:310:28
        rob_uop_20_edge_inst = _RANDOM[11'h117][24];	// rob.scala:310:28
        rob_uop_20_pc_lob = _RANDOM[11'h117][30:25];	// rob.scala:310:28
        rob_uop_20_pdst = _RANDOM[11'h119][25:19];	// rob.scala:310:28
        rob_uop_20_stale_pdst = _RANDOM[11'h11A][30:24];	// rob.scala:310:28
        rob_uop_20_is_fencei = _RANDOM[11'h11D][10];	// rob.scala:310:28
        rob_uop_20_uses_ldq = _RANDOM[11'h11D][12];	// rob.scala:310:28
        rob_uop_20_uses_stq = _RANDOM[11'h11D][13];	// rob.scala:310:28
        rob_uop_20_is_sys_pc2epc = _RANDOM[11'h11D][14];	// rob.scala:310:28
        rob_uop_20_flush_on_commit = _RANDOM[11'h11D][16];	// rob.scala:310:28
        rob_uop_20_ldst = _RANDOM[11'h11D][23:18];	// rob.scala:310:28
        rob_uop_20_ldst_val = _RANDOM[11'h11E][10];	// rob.scala:310:28
        rob_uop_20_dst_rtype = _RANDOM[11'h11E][12:11];	// rob.scala:310:28
        rob_uop_20_fp_val = _RANDOM[11'h11E][18];	// rob.scala:310:28
        rob_uop_21_uopc = {_RANDOM[11'h11E][31:29], _RANDOM[11'h11F][3:0]};	// rob.scala:310:28
        rob_uop_21_is_rvc = _RANDOM[11'h121][4];	// rob.scala:310:28
        rob_uop_21_br_mask = {_RANDOM[11'h123][31:25], _RANDOM[11'h124][8:0]};	// rob.scala:310:28
        rob_uop_21_ftq_idx = _RANDOM[11'h124][17:13];	// rob.scala:310:28
        rob_uop_21_edge_inst = _RANDOM[11'h124][18];	// rob.scala:310:28
        rob_uop_21_pc_lob = _RANDOM[11'h124][24:19];	// rob.scala:310:28
        rob_uop_21_pdst = _RANDOM[11'h126][19:13];	// rob.scala:310:28
        rob_uop_21_stale_pdst = _RANDOM[11'h127][24:18];	// rob.scala:310:28
        rob_uop_21_is_fencei = _RANDOM[11'h12A][4];	// rob.scala:310:28
        rob_uop_21_uses_ldq = _RANDOM[11'h12A][6];	// rob.scala:310:28
        rob_uop_21_uses_stq = _RANDOM[11'h12A][7];	// rob.scala:310:28
        rob_uop_21_is_sys_pc2epc = _RANDOM[11'h12A][8];	// rob.scala:310:28
        rob_uop_21_flush_on_commit = _RANDOM[11'h12A][10];	// rob.scala:310:28
        rob_uop_21_ldst = _RANDOM[11'h12A][17:12];	// rob.scala:310:28
        rob_uop_21_ldst_val = _RANDOM[11'h12B][4];	// rob.scala:310:28
        rob_uop_21_dst_rtype = _RANDOM[11'h12B][6:5];	// rob.scala:310:28
        rob_uop_21_fp_val = _RANDOM[11'h12B][12];	// rob.scala:310:28
        rob_uop_22_uopc = _RANDOM[11'h12B][29:23];	// rob.scala:310:28
        rob_uop_22_is_rvc = _RANDOM[11'h12D][30];	// rob.scala:310:28
        rob_uop_22_br_mask = {_RANDOM[11'h130][31:19], _RANDOM[11'h131][2:0]};	// rob.scala:310:28
        rob_uop_22_ftq_idx = _RANDOM[11'h131][11:7];	// rob.scala:310:28
        rob_uop_22_edge_inst = _RANDOM[11'h131][12];	// rob.scala:310:28
        rob_uop_22_pc_lob = _RANDOM[11'h131][18:13];	// rob.scala:310:28
        rob_uop_22_pdst = _RANDOM[11'h133][13:7];	// rob.scala:310:28
        rob_uop_22_stale_pdst = _RANDOM[11'h134][18:12];	// rob.scala:310:28
        rob_uop_22_is_fencei = _RANDOM[11'h136][30];	// rob.scala:310:28
        rob_uop_22_uses_ldq = _RANDOM[11'h137][0];	// rob.scala:310:28
        rob_uop_22_uses_stq = _RANDOM[11'h137][1];	// rob.scala:310:28
        rob_uop_22_is_sys_pc2epc = _RANDOM[11'h137][2];	// rob.scala:310:28
        rob_uop_22_flush_on_commit = _RANDOM[11'h137][4];	// rob.scala:310:28
        rob_uop_22_ldst = _RANDOM[11'h137][11:6];	// rob.scala:310:28
        rob_uop_22_ldst_val = _RANDOM[11'h137][30];	// rob.scala:310:28
        rob_uop_22_dst_rtype = {_RANDOM[11'h137][31], _RANDOM[11'h138][0]};	// rob.scala:310:28
        rob_uop_22_fp_val = _RANDOM[11'h138][6];	// rob.scala:310:28
        rob_uop_23_uopc = _RANDOM[11'h138][23:17];	// rob.scala:310:28
        rob_uop_23_is_rvc = _RANDOM[11'h13A][24];	// rob.scala:310:28
        rob_uop_23_br_mask = _RANDOM[11'h13D][28:13];	// rob.scala:310:28
        rob_uop_23_ftq_idx = _RANDOM[11'h13E][5:1];	// rob.scala:310:28
        rob_uop_23_edge_inst = _RANDOM[11'h13E][6];	// rob.scala:310:28
        rob_uop_23_pc_lob = _RANDOM[11'h13E][12:7];	// rob.scala:310:28
        rob_uop_23_pdst = _RANDOM[11'h140][7:1];	// rob.scala:310:28
        rob_uop_23_stale_pdst = _RANDOM[11'h141][12:6];	// rob.scala:310:28
        rob_uop_23_is_fencei = _RANDOM[11'h143][24];	// rob.scala:310:28
        rob_uop_23_uses_ldq = _RANDOM[11'h143][26];	// rob.scala:310:28
        rob_uop_23_uses_stq = _RANDOM[11'h143][27];	// rob.scala:310:28
        rob_uop_23_is_sys_pc2epc = _RANDOM[11'h143][28];	// rob.scala:310:28
        rob_uop_23_flush_on_commit = _RANDOM[11'h143][30];	// rob.scala:310:28
        rob_uop_23_ldst = _RANDOM[11'h144][5:0];	// rob.scala:310:28
        rob_uop_23_ldst_val = _RANDOM[11'h144][24];	// rob.scala:310:28
        rob_uop_23_dst_rtype = _RANDOM[11'h144][26:25];	// rob.scala:310:28
        rob_uop_23_fp_val = _RANDOM[11'h145][0];	// rob.scala:310:28
        rob_uop_24_uopc = _RANDOM[11'h145][17:11];	// rob.scala:310:28
        rob_uop_24_is_rvc = _RANDOM[11'h147][18];	// rob.scala:310:28
        rob_uop_24_br_mask = _RANDOM[11'h14A][22:7];	// rob.scala:310:28
        rob_uop_24_ftq_idx = _RANDOM[11'h14A][31:27];	// rob.scala:310:28
        rob_uop_24_edge_inst = _RANDOM[11'h14B][0];	// rob.scala:310:28
        rob_uop_24_pc_lob = _RANDOM[11'h14B][6:1];	// rob.scala:310:28
        rob_uop_24_pdst = {_RANDOM[11'h14C][31:27], _RANDOM[11'h14D][1:0]};	// rob.scala:310:28
        rob_uop_24_stale_pdst = _RANDOM[11'h14E][6:0];	// rob.scala:310:28
        rob_uop_24_is_fencei = _RANDOM[11'h150][18];	// rob.scala:310:28
        rob_uop_24_uses_ldq = _RANDOM[11'h150][20];	// rob.scala:310:28
        rob_uop_24_uses_stq = _RANDOM[11'h150][21];	// rob.scala:310:28
        rob_uop_24_is_sys_pc2epc = _RANDOM[11'h150][22];	// rob.scala:310:28
        rob_uop_24_flush_on_commit = _RANDOM[11'h150][24];	// rob.scala:310:28
        rob_uop_24_ldst = _RANDOM[11'h150][31:26];	// rob.scala:310:28
        rob_uop_24_ldst_val = _RANDOM[11'h151][18];	// rob.scala:310:28
        rob_uop_24_dst_rtype = _RANDOM[11'h151][20:19];	// rob.scala:310:28
        rob_uop_24_fp_val = _RANDOM[11'h151][26];	// rob.scala:310:28
        rob_uop_25_uopc = _RANDOM[11'h152][11:5];	// rob.scala:310:28
        rob_uop_25_is_rvc = _RANDOM[11'h154][12];	// rob.scala:310:28
        rob_uop_25_br_mask = _RANDOM[11'h157][16:1];	// rob.scala:310:28
        rob_uop_25_ftq_idx = _RANDOM[11'h157][25:21];	// rob.scala:310:28
        rob_uop_25_edge_inst = _RANDOM[11'h157][26];	// rob.scala:310:28
        rob_uop_25_pc_lob = {_RANDOM[11'h157][31:27], _RANDOM[11'h158][0]};	// rob.scala:310:28
        rob_uop_25_pdst = _RANDOM[11'h159][27:21];	// rob.scala:310:28
        rob_uop_25_stale_pdst = {_RANDOM[11'h15A][31:26], _RANDOM[11'h15B][0]};	// rob.scala:310:28
        rob_uop_25_is_fencei = _RANDOM[11'h15D][12];	// rob.scala:310:28
        rob_uop_25_uses_ldq = _RANDOM[11'h15D][14];	// rob.scala:310:28
        rob_uop_25_uses_stq = _RANDOM[11'h15D][15];	// rob.scala:310:28
        rob_uop_25_is_sys_pc2epc = _RANDOM[11'h15D][16];	// rob.scala:310:28
        rob_uop_25_flush_on_commit = _RANDOM[11'h15D][18];	// rob.scala:310:28
        rob_uop_25_ldst = _RANDOM[11'h15D][25:20];	// rob.scala:310:28
        rob_uop_25_ldst_val = _RANDOM[11'h15E][12];	// rob.scala:310:28
        rob_uop_25_dst_rtype = _RANDOM[11'h15E][14:13];	// rob.scala:310:28
        rob_uop_25_fp_val = _RANDOM[11'h15E][20];	// rob.scala:310:28
        rob_uop_26_uopc = {_RANDOM[11'h15E][31], _RANDOM[11'h15F][5:0]};	// rob.scala:310:28
        rob_uop_26_is_rvc = _RANDOM[11'h161][6];	// rob.scala:310:28
        rob_uop_26_br_mask = {_RANDOM[11'h163][31:27], _RANDOM[11'h164][10:0]};	// rob.scala:310:28
        rob_uop_26_ftq_idx = _RANDOM[11'h164][19:15];	// rob.scala:310:28
        rob_uop_26_edge_inst = _RANDOM[11'h164][20];	// rob.scala:310:28
        rob_uop_26_pc_lob = _RANDOM[11'h164][26:21];	// rob.scala:310:28
        rob_uop_26_pdst = _RANDOM[11'h166][21:15];	// rob.scala:310:28
        rob_uop_26_stale_pdst = _RANDOM[11'h167][26:20];	// rob.scala:310:28
        rob_uop_26_is_fencei = _RANDOM[11'h16A][6];	// rob.scala:310:28
        rob_uop_26_uses_ldq = _RANDOM[11'h16A][8];	// rob.scala:310:28
        rob_uop_26_uses_stq = _RANDOM[11'h16A][9];	// rob.scala:310:28
        rob_uop_26_is_sys_pc2epc = _RANDOM[11'h16A][10];	// rob.scala:310:28
        rob_uop_26_flush_on_commit = _RANDOM[11'h16A][12];	// rob.scala:310:28
        rob_uop_26_ldst = _RANDOM[11'h16A][19:14];	// rob.scala:310:28
        rob_uop_26_ldst_val = _RANDOM[11'h16B][6];	// rob.scala:310:28
        rob_uop_26_dst_rtype = _RANDOM[11'h16B][8:7];	// rob.scala:310:28
        rob_uop_26_fp_val = _RANDOM[11'h16B][14];	// rob.scala:310:28
        rob_uop_27_uopc = _RANDOM[11'h16B][31:25];	// rob.scala:310:28
        rob_uop_27_is_rvc = _RANDOM[11'h16E][0];	// rob.scala:310:28
        rob_uop_27_br_mask = {_RANDOM[11'h170][31:21], _RANDOM[11'h171][4:0]};	// rob.scala:310:28
        rob_uop_27_ftq_idx = _RANDOM[11'h171][13:9];	// rob.scala:310:28
        rob_uop_27_edge_inst = _RANDOM[11'h171][14];	// rob.scala:310:28
        rob_uop_27_pc_lob = _RANDOM[11'h171][20:15];	// rob.scala:310:28
        rob_uop_27_pdst = _RANDOM[11'h173][15:9];	// rob.scala:310:28
        rob_uop_27_stale_pdst = _RANDOM[11'h174][20:14];	// rob.scala:310:28
        rob_uop_27_is_fencei = _RANDOM[11'h177][0];	// rob.scala:310:28
        rob_uop_27_uses_ldq = _RANDOM[11'h177][2];	// rob.scala:310:28
        rob_uop_27_uses_stq = _RANDOM[11'h177][3];	// rob.scala:310:28
        rob_uop_27_is_sys_pc2epc = _RANDOM[11'h177][4];	// rob.scala:310:28
        rob_uop_27_flush_on_commit = _RANDOM[11'h177][6];	// rob.scala:310:28
        rob_uop_27_ldst = _RANDOM[11'h177][13:8];	// rob.scala:310:28
        rob_uop_27_ldst_val = _RANDOM[11'h178][0];	// rob.scala:310:28
        rob_uop_27_dst_rtype = _RANDOM[11'h178][2:1];	// rob.scala:310:28
        rob_uop_27_fp_val = _RANDOM[11'h178][8];	// rob.scala:310:28
        rob_uop_28_uopc = _RANDOM[11'h178][25:19];	// rob.scala:310:28
        rob_uop_28_is_rvc = _RANDOM[11'h17A][26];	// rob.scala:310:28
        rob_uop_28_br_mask = _RANDOM[11'h17D][30:15];	// rob.scala:310:28
        rob_uop_28_ftq_idx = _RANDOM[11'h17E][7:3];	// rob.scala:310:28
        rob_uop_28_edge_inst = _RANDOM[11'h17E][8];	// rob.scala:310:28
        rob_uop_28_pc_lob = _RANDOM[11'h17E][14:9];	// rob.scala:310:28
        rob_uop_28_pdst = _RANDOM[11'h180][9:3];	// rob.scala:310:28
        rob_uop_28_stale_pdst = _RANDOM[11'h181][14:8];	// rob.scala:310:28
        rob_uop_28_is_fencei = _RANDOM[11'h183][26];	// rob.scala:310:28
        rob_uop_28_uses_ldq = _RANDOM[11'h183][28];	// rob.scala:310:28
        rob_uop_28_uses_stq = _RANDOM[11'h183][29];	// rob.scala:310:28
        rob_uop_28_is_sys_pc2epc = _RANDOM[11'h183][30];	// rob.scala:310:28
        rob_uop_28_flush_on_commit = _RANDOM[11'h184][0];	// rob.scala:310:28
        rob_uop_28_ldst = _RANDOM[11'h184][7:2];	// rob.scala:310:28
        rob_uop_28_ldst_val = _RANDOM[11'h184][26];	// rob.scala:310:28
        rob_uop_28_dst_rtype = _RANDOM[11'h184][28:27];	// rob.scala:310:28
        rob_uop_28_fp_val = _RANDOM[11'h185][2];	// rob.scala:310:28
        rob_uop_29_uopc = _RANDOM[11'h185][19:13];	// rob.scala:310:28
        rob_uop_29_is_rvc = _RANDOM[11'h187][20];	// rob.scala:310:28
        rob_uop_29_br_mask = _RANDOM[11'h18A][24:9];	// rob.scala:310:28
        rob_uop_29_ftq_idx = {_RANDOM[11'h18A][31:29], _RANDOM[11'h18B][1:0]};	// rob.scala:310:28
        rob_uop_29_edge_inst = _RANDOM[11'h18B][2];	// rob.scala:310:28
        rob_uop_29_pc_lob = _RANDOM[11'h18B][8:3];	// rob.scala:310:28
        rob_uop_29_pdst = {_RANDOM[11'h18C][31:29], _RANDOM[11'h18D][3:0]};	// rob.scala:310:28
        rob_uop_29_stale_pdst = _RANDOM[11'h18E][8:2];	// rob.scala:310:28
        rob_uop_29_is_fencei = _RANDOM[11'h190][20];	// rob.scala:310:28
        rob_uop_29_uses_ldq = _RANDOM[11'h190][22];	// rob.scala:310:28
        rob_uop_29_uses_stq = _RANDOM[11'h190][23];	// rob.scala:310:28
        rob_uop_29_is_sys_pc2epc = _RANDOM[11'h190][24];	// rob.scala:310:28
        rob_uop_29_flush_on_commit = _RANDOM[11'h190][26];	// rob.scala:310:28
        rob_uop_29_ldst = {_RANDOM[11'h190][31:28], _RANDOM[11'h191][1:0]};	// rob.scala:310:28
        rob_uop_29_ldst_val = _RANDOM[11'h191][20];	// rob.scala:310:28
        rob_uop_29_dst_rtype = _RANDOM[11'h191][22:21];	// rob.scala:310:28
        rob_uop_29_fp_val = _RANDOM[11'h191][28];	// rob.scala:310:28
        rob_uop_30_uopc = _RANDOM[11'h192][13:7];	// rob.scala:310:28
        rob_uop_30_is_rvc = _RANDOM[11'h194][14];	// rob.scala:310:28
        rob_uop_30_br_mask = _RANDOM[11'h197][18:3];	// rob.scala:310:28
        rob_uop_30_ftq_idx = _RANDOM[11'h197][27:23];	// rob.scala:310:28
        rob_uop_30_edge_inst = _RANDOM[11'h197][28];	// rob.scala:310:28
        rob_uop_30_pc_lob = {_RANDOM[11'h197][31:29], _RANDOM[11'h198][2:0]};	// rob.scala:310:28
        rob_uop_30_pdst = _RANDOM[11'h199][29:23];	// rob.scala:310:28
        rob_uop_30_stale_pdst = {_RANDOM[11'h19A][31:28], _RANDOM[11'h19B][2:0]};	// rob.scala:310:28
        rob_uop_30_is_fencei = _RANDOM[11'h19D][14];	// rob.scala:310:28
        rob_uop_30_uses_ldq = _RANDOM[11'h19D][16];	// rob.scala:310:28
        rob_uop_30_uses_stq = _RANDOM[11'h19D][17];	// rob.scala:310:28
        rob_uop_30_is_sys_pc2epc = _RANDOM[11'h19D][18];	// rob.scala:310:28
        rob_uop_30_flush_on_commit = _RANDOM[11'h19D][20];	// rob.scala:310:28
        rob_uop_30_ldst = _RANDOM[11'h19D][27:22];	// rob.scala:310:28
        rob_uop_30_ldst_val = _RANDOM[11'h19E][14];	// rob.scala:310:28
        rob_uop_30_dst_rtype = _RANDOM[11'h19E][16:15];	// rob.scala:310:28
        rob_uop_30_fp_val = _RANDOM[11'h19E][22];	// rob.scala:310:28
        rob_uop_31_uopc = _RANDOM[11'h19F][7:1];	// rob.scala:310:28
        rob_uop_31_is_rvc = _RANDOM[11'h1A1][8];	// rob.scala:310:28
        rob_uop_31_br_mask = {_RANDOM[11'h1A3][31:29], _RANDOM[11'h1A4][12:0]};	// rob.scala:310:28
        rob_uop_31_ftq_idx = _RANDOM[11'h1A4][21:17];	// rob.scala:310:28
        rob_uop_31_edge_inst = _RANDOM[11'h1A4][22];	// rob.scala:310:28
        rob_uop_31_pc_lob = _RANDOM[11'h1A4][28:23];	// rob.scala:310:28
        rob_uop_31_pdst = _RANDOM[11'h1A6][23:17];	// rob.scala:310:28
        rob_uop_31_stale_pdst = _RANDOM[11'h1A7][28:22];	// rob.scala:310:28
        rob_uop_31_is_fencei = _RANDOM[11'h1AA][8];	// rob.scala:310:28
        rob_uop_31_uses_ldq = _RANDOM[11'h1AA][10];	// rob.scala:310:28
        rob_uop_31_uses_stq = _RANDOM[11'h1AA][11];	// rob.scala:310:28
        rob_uop_31_is_sys_pc2epc = _RANDOM[11'h1AA][12];	// rob.scala:310:28
        rob_uop_31_flush_on_commit = _RANDOM[11'h1AA][14];	// rob.scala:310:28
        rob_uop_31_ldst = _RANDOM[11'h1AA][21:16];	// rob.scala:310:28
        rob_uop_31_ldst_val = _RANDOM[11'h1AB][8];	// rob.scala:310:28
        rob_uop_31_dst_rtype = _RANDOM[11'h1AB][10:9];	// rob.scala:310:28
        rob_uop_31_fp_val = _RANDOM[11'h1AB][16];	// rob.scala:310:28
        rob_exception_0 = _RANDOM[11'h1AB][27];	// rob.scala:310:28, :311:28
        rob_exception_1 = _RANDOM[11'h1AB][28];	// rob.scala:310:28, :311:28
        rob_exception_2 = _RANDOM[11'h1AB][29];	// rob.scala:310:28, :311:28
        rob_exception_3 = _RANDOM[11'h1AB][30];	// rob.scala:310:28, :311:28
        rob_exception_4 = _RANDOM[11'h1AB][31];	// rob.scala:310:28, :311:28
        rob_exception_5 = _RANDOM[11'h1AC][0];	// rob.scala:311:28
        rob_exception_6 = _RANDOM[11'h1AC][1];	// rob.scala:311:28
        rob_exception_7 = _RANDOM[11'h1AC][2];	// rob.scala:311:28
        rob_exception_8 = _RANDOM[11'h1AC][3];	// rob.scala:311:28
        rob_exception_9 = _RANDOM[11'h1AC][4];	// rob.scala:311:28
        rob_exception_10 = _RANDOM[11'h1AC][5];	// rob.scala:311:28
        rob_exception_11 = _RANDOM[11'h1AC][6];	// rob.scala:311:28
        rob_exception_12 = _RANDOM[11'h1AC][7];	// rob.scala:311:28
        rob_exception_13 = _RANDOM[11'h1AC][8];	// rob.scala:311:28
        rob_exception_14 = _RANDOM[11'h1AC][9];	// rob.scala:311:28
        rob_exception_15 = _RANDOM[11'h1AC][10];	// rob.scala:311:28
        rob_exception_16 = _RANDOM[11'h1AC][11];	// rob.scala:311:28
        rob_exception_17 = _RANDOM[11'h1AC][12];	// rob.scala:311:28
        rob_exception_18 = _RANDOM[11'h1AC][13];	// rob.scala:311:28
        rob_exception_19 = _RANDOM[11'h1AC][14];	// rob.scala:311:28
        rob_exception_20 = _RANDOM[11'h1AC][15];	// rob.scala:311:28
        rob_exception_21 = _RANDOM[11'h1AC][16];	// rob.scala:311:28
        rob_exception_22 = _RANDOM[11'h1AC][17];	// rob.scala:311:28
        rob_exception_23 = _RANDOM[11'h1AC][18];	// rob.scala:311:28
        rob_exception_24 = _RANDOM[11'h1AC][19];	// rob.scala:311:28
        rob_exception_25 = _RANDOM[11'h1AC][20];	// rob.scala:311:28
        rob_exception_26 = _RANDOM[11'h1AC][21];	// rob.scala:311:28
        rob_exception_27 = _RANDOM[11'h1AC][22];	// rob.scala:311:28
        rob_exception_28 = _RANDOM[11'h1AC][23];	// rob.scala:311:28
        rob_exception_29 = _RANDOM[11'h1AC][24];	// rob.scala:311:28
        rob_exception_30 = _RANDOM[11'h1AC][25];	// rob.scala:311:28
        rob_exception_31 = _RANDOM[11'h1AC][26];	// rob.scala:311:28
        rob_predicated_0 = _RANDOM[11'h1AC][27];	// rob.scala:311:28, :312:29
        rob_predicated_1 = _RANDOM[11'h1AC][28];	// rob.scala:311:28, :312:29
        rob_predicated_2 = _RANDOM[11'h1AC][29];	// rob.scala:311:28, :312:29
        rob_predicated_3 = _RANDOM[11'h1AC][30];	// rob.scala:311:28, :312:29
        rob_predicated_4 = _RANDOM[11'h1AC][31];	// rob.scala:311:28, :312:29
        rob_predicated_5 = _RANDOM[11'h1AD][0];	// rob.scala:312:29
        rob_predicated_6 = _RANDOM[11'h1AD][1];	// rob.scala:312:29
        rob_predicated_7 = _RANDOM[11'h1AD][2];	// rob.scala:312:29
        rob_predicated_8 = _RANDOM[11'h1AD][3];	// rob.scala:312:29
        rob_predicated_9 = _RANDOM[11'h1AD][4];	// rob.scala:312:29
        rob_predicated_10 = _RANDOM[11'h1AD][5];	// rob.scala:312:29
        rob_predicated_11 = _RANDOM[11'h1AD][6];	// rob.scala:312:29
        rob_predicated_12 = _RANDOM[11'h1AD][7];	// rob.scala:312:29
        rob_predicated_13 = _RANDOM[11'h1AD][8];	// rob.scala:312:29
        rob_predicated_14 = _RANDOM[11'h1AD][9];	// rob.scala:312:29
        rob_predicated_15 = _RANDOM[11'h1AD][10];	// rob.scala:312:29
        rob_predicated_16 = _RANDOM[11'h1AD][11];	// rob.scala:312:29
        rob_predicated_17 = _RANDOM[11'h1AD][12];	// rob.scala:312:29
        rob_predicated_18 = _RANDOM[11'h1AD][13];	// rob.scala:312:29
        rob_predicated_19 = _RANDOM[11'h1AD][14];	// rob.scala:312:29
        rob_predicated_20 = _RANDOM[11'h1AD][15];	// rob.scala:312:29
        rob_predicated_21 = _RANDOM[11'h1AD][16];	// rob.scala:312:29
        rob_predicated_22 = _RANDOM[11'h1AD][17];	// rob.scala:312:29
        rob_predicated_23 = _RANDOM[11'h1AD][18];	// rob.scala:312:29
        rob_predicated_24 = _RANDOM[11'h1AD][19];	// rob.scala:312:29
        rob_predicated_25 = _RANDOM[11'h1AD][20];	// rob.scala:312:29
        rob_predicated_26 = _RANDOM[11'h1AD][21];	// rob.scala:312:29
        rob_predicated_27 = _RANDOM[11'h1AD][22];	// rob.scala:312:29
        rob_predicated_28 = _RANDOM[11'h1AD][23];	// rob.scala:312:29
        rob_predicated_29 = _RANDOM[11'h1AD][24];	// rob.scala:312:29
        rob_predicated_30 = _RANDOM[11'h1AD][25];	// rob.scala:312:29
        rob_predicated_31 = _RANDOM[11'h1AD][26];	// rob.scala:312:29
        rob_val_1_0 = _RANDOM[11'h1AD][27];	// rob.scala:307:32, :312:29
        rob_val_1_1 = _RANDOM[11'h1AD][28];	// rob.scala:307:32, :312:29
        rob_val_1_2 = _RANDOM[11'h1AD][29];	// rob.scala:307:32, :312:29
        rob_val_1_3 = _RANDOM[11'h1AD][30];	// rob.scala:307:32, :312:29
        rob_val_1_4 = _RANDOM[11'h1AD][31];	// rob.scala:307:32, :312:29
        rob_val_1_5 = _RANDOM[11'h1AE][0];	// rob.scala:307:32
        rob_val_1_6 = _RANDOM[11'h1AE][1];	// rob.scala:307:32
        rob_val_1_7 = _RANDOM[11'h1AE][2];	// rob.scala:307:32
        rob_val_1_8 = _RANDOM[11'h1AE][3];	// rob.scala:307:32
        rob_val_1_9 = _RANDOM[11'h1AE][4];	// rob.scala:307:32
        rob_val_1_10 = _RANDOM[11'h1AE][5];	// rob.scala:307:32
        rob_val_1_11 = _RANDOM[11'h1AE][6];	// rob.scala:307:32
        rob_val_1_12 = _RANDOM[11'h1AE][7];	// rob.scala:307:32
        rob_val_1_13 = _RANDOM[11'h1AE][8];	// rob.scala:307:32
        rob_val_1_14 = _RANDOM[11'h1AE][9];	// rob.scala:307:32
        rob_val_1_15 = _RANDOM[11'h1AE][10];	// rob.scala:307:32
        rob_val_1_16 = _RANDOM[11'h1AE][11];	// rob.scala:307:32
        rob_val_1_17 = _RANDOM[11'h1AE][12];	// rob.scala:307:32
        rob_val_1_18 = _RANDOM[11'h1AE][13];	// rob.scala:307:32
        rob_val_1_19 = _RANDOM[11'h1AE][14];	// rob.scala:307:32
        rob_val_1_20 = _RANDOM[11'h1AE][15];	// rob.scala:307:32
        rob_val_1_21 = _RANDOM[11'h1AE][16];	// rob.scala:307:32
        rob_val_1_22 = _RANDOM[11'h1AE][17];	// rob.scala:307:32
        rob_val_1_23 = _RANDOM[11'h1AE][18];	// rob.scala:307:32
        rob_val_1_24 = _RANDOM[11'h1AE][19];	// rob.scala:307:32
        rob_val_1_25 = _RANDOM[11'h1AE][20];	// rob.scala:307:32
        rob_val_1_26 = _RANDOM[11'h1AE][21];	// rob.scala:307:32
        rob_val_1_27 = _RANDOM[11'h1AE][22];	// rob.scala:307:32
        rob_val_1_28 = _RANDOM[11'h1AE][23];	// rob.scala:307:32
        rob_val_1_29 = _RANDOM[11'h1AE][24];	// rob.scala:307:32
        rob_val_1_30 = _RANDOM[11'h1AE][25];	// rob.scala:307:32
        rob_val_1_31 = _RANDOM[11'h1AE][26];	// rob.scala:307:32
        rob_bsy_1_0 = _RANDOM[11'h1AE][27];	// rob.scala:307:32, :308:28
        rob_bsy_1_1 = _RANDOM[11'h1AE][28];	// rob.scala:307:32, :308:28
        rob_bsy_1_2 = _RANDOM[11'h1AE][29];	// rob.scala:307:32, :308:28
        rob_bsy_1_3 = _RANDOM[11'h1AE][30];	// rob.scala:307:32, :308:28
        rob_bsy_1_4 = _RANDOM[11'h1AE][31];	// rob.scala:307:32, :308:28
        rob_bsy_1_5 = _RANDOM[11'h1AF][0];	// rob.scala:308:28
        rob_bsy_1_6 = _RANDOM[11'h1AF][1];	// rob.scala:308:28
        rob_bsy_1_7 = _RANDOM[11'h1AF][2];	// rob.scala:308:28
        rob_bsy_1_8 = _RANDOM[11'h1AF][3];	// rob.scala:308:28
        rob_bsy_1_9 = _RANDOM[11'h1AF][4];	// rob.scala:308:28
        rob_bsy_1_10 = _RANDOM[11'h1AF][5];	// rob.scala:308:28
        rob_bsy_1_11 = _RANDOM[11'h1AF][6];	// rob.scala:308:28
        rob_bsy_1_12 = _RANDOM[11'h1AF][7];	// rob.scala:308:28
        rob_bsy_1_13 = _RANDOM[11'h1AF][8];	// rob.scala:308:28
        rob_bsy_1_14 = _RANDOM[11'h1AF][9];	// rob.scala:308:28
        rob_bsy_1_15 = _RANDOM[11'h1AF][10];	// rob.scala:308:28
        rob_bsy_1_16 = _RANDOM[11'h1AF][11];	// rob.scala:308:28
        rob_bsy_1_17 = _RANDOM[11'h1AF][12];	// rob.scala:308:28
        rob_bsy_1_18 = _RANDOM[11'h1AF][13];	// rob.scala:308:28
        rob_bsy_1_19 = _RANDOM[11'h1AF][14];	// rob.scala:308:28
        rob_bsy_1_20 = _RANDOM[11'h1AF][15];	// rob.scala:308:28
        rob_bsy_1_21 = _RANDOM[11'h1AF][16];	// rob.scala:308:28
        rob_bsy_1_22 = _RANDOM[11'h1AF][17];	// rob.scala:308:28
        rob_bsy_1_23 = _RANDOM[11'h1AF][18];	// rob.scala:308:28
        rob_bsy_1_24 = _RANDOM[11'h1AF][19];	// rob.scala:308:28
        rob_bsy_1_25 = _RANDOM[11'h1AF][20];	// rob.scala:308:28
        rob_bsy_1_26 = _RANDOM[11'h1AF][21];	// rob.scala:308:28
        rob_bsy_1_27 = _RANDOM[11'h1AF][22];	// rob.scala:308:28
        rob_bsy_1_28 = _RANDOM[11'h1AF][23];	// rob.scala:308:28
        rob_bsy_1_29 = _RANDOM[11'h1AF][24];	// rob.scala:308:28
        rob_bsy_1_30 = _RANDOM[11'h1AF][25];	// rob.scala:308:28
        rob_bsy_1_31 = _RANDOM[11'h1AF][26];	// rob.scala:308:28
        rob_unsafe_1_0 = _RANDOM[11'h1AF][27];	// rob.scala:308:28, :309:28
        rob_unsafe_1_1 = _RANDOM[11'h1AF][28];	// rob.scala:308:28, :309:28
        rob_unsafe_1_2 = _RANDOM[11'h1AF][29];	// rob.scala:308:28, :309:28
        rob_unsafe_1_3 = _RANDOM[11'h1AF][30];	// rob.scala:308:28, :309:28
        rob_unsafe_1_4 = _RANDOM[11'h1AF][31];	// rob.scala:308:28, :309:28
        rob_unsafe_1_5 = _RANDOM[11'h1B0][0];	// rob.scala:309:28
        rob_unsafe_1_6 = _RANDOM[11'h1B0][1];	// rob.scala:309:28
        rob_unsafe_1_7 = _RANDOM[11'h1B0][2];	// rob.scala:309:28
        rob_unsafe_1_8 = _RANDOM[11'h1B0][3];	// rob.scala:309:28
        rob_unsafe_1_9 = _RANDOM[11'h1B0][4];	// rob.scala:309:28
        rob_unsafe_1_10 = _RANDOM[11'h1B0][5];	// rob.scala:309:28
        rob_unsafe_1_11 = _RANDOM[11'h1B0][6];	// rob.scala:309:28
        rob_unsafe_1_12 = _RANDOM[11'h1B0][7];	// rob.scala:309:28
        rob_unsafe_1_13 = _RANDOM[11'h1B0][8];	// rob.scala:309:28
        rob_unsafe_1_14 = _RANDOM[11'h1B0][9];	// rob.scala:309:28
        rob_unsafe_1_15 = _RANDOM[11'h1B0][10];	// rob.scala:309:28
        rob_unsafe_1_16 = _RANDOM[11'h1B0][11];	// rob.scala:309:28
        rob_unsafe_1_17 = _RANDOM[11'h1B0][12];	// rob.scala:309:28
        rob_unsafe_1_18 = _RANDOM[11'h1B0][13];	// rob.scala:309:28
        rob_unsafe_1_19 = _RANDOM[11'h1B0][14];	// rob.scala:309:28
        rob_unsafe_1_20 = _RANDOM[11'h1B0][15];	// rob.scala:309:28
        rob_unsafe_1_21 = _RANDOM[11'h1B0][16];	// rob.scala:309:28
        rob_unsafe_1_22 = _RANDOM[11'h1B0][17];	// rob.scala:309:28
        rob_unsafe_1_23 = _RANDOM[11'h1B0][18];	// rob.scala:309:28
        rob_unsafe_1_24 = _RANDOM[11'h1B0][19];	// rob.scala:309:28
        rob_unsafe_1_25 = _RANDOM[11'h1B0][20];	// rob.scala:309:28
        rob_unsafe_1_26 = _RANDOM[11'h1B0][21];	// rob.scala:309:28
        rob_unsafe_1_27 = _RANDOM[11'h1B0][22];	// rob.scala:309:28
        rob_unsafe_1_28 = _RANDOM[11'h1B0][23];	// rob.scala:309:28
        rob_unsafe_1_29 = _RANDOM[11'h1B0][24];	// rob.scala:309:28
        rob_unsafe_1_30 = _RANDOM[11'h1B0][25];	// rob.scala:309:28
        rob_unsafe_1_31 = _RANDOM[11'h1B0][26];	// rob.scala:309:28
        rob_uop_1_0_uopc = {_RANDOM[11'h1B0][31:27], _RANDOM[11'h1B1][1:0]};	// rob.scala:309:28, :310:28
        rob_uop_1_0_is_rvc = _RANDOM[11'h1B3][2];	// rob.scala:310:28
        rob_uop_1_0_br_mask = {_RANDOM[11'h1B5][31:23], _RANDOM[11'h1B6][6:0]};	// rob.scala:310:28
        rob_uop_1_0_ftq_idx = _RANDOM[11'h1B6][15:11];	// rob.scala:310:28
        rob_uop_1_0_edge_inst = _RANDOM[11'h1B6][16];	// rob.scala:310:28
        rob_uop_1_0_pc_lob = _RANDOM[11'h1B6][22:17];	// rob.scala:310:28
        rob_uop_1_0_pdst = _RANDOM[11'h1B8][17:11];	// rob.scala:310:28
        rob_uop_1_0_stale_pdst = _RANDOM[11'h1B9][22:16];	// rob.scala:310:28
        rob_uop_1_0_is_fencei = _RANDOM[11'h1BC][2];	// rob.scala:310:28
        rob_uop_1_0_uses_ldq = _RANDOM[11'h1BC][4];	// rob.scala:310:28
        rob_uop_1_0_uses_stq = _RANDOM[11'h1BC][5];	// rob.scala:310:28
        rob_uop_1_0_is_sys_pc2epc = _RANDOM[11'h1BC][6];	// rob.scala:310:28
        rob_uop_1_0_flush_on_commit = _RANDOM[11'h1BC][8];	// rob.scala:310:28
        rob_uop_1_0_ldst = _RANDOM[11'h1BC][15:10];	// rob.scala:310:28
        rob_uop_1_0_ldst_val = _RANDOM[11'h1BD][2];	// rob.scala:310:28
        rob_uop_1_0_dst_rtype = _RANDOM[11'h1BD][4:3];	// rob.scala:310:28
        rob_uop_1_0_fp_val = _RANDOM[11'h1BD][10];	// rob.scala:310:28
        rob_uop_1_1_uopc = _RANDOM[11'h1BD][27:21];	// rob.scala:310:28
        rob_uop_1_1_is_rvc = _RANDOM[11'h1BF][28];	// rob.scala:310:28
        rob_uop_1_1_br_mask = {_RANDOM[11'h1C2][31:17], _RANDOM[11'h1C3][0]};	// rob.scala:310:28
        rob_uop_1_1_ftq_idx = _RANDOM[11'h1C3][9:5];	// rob.scala:310:28
        rob_uop_1_1_edge_inst = _RANDOM[11'h1C3][10];	// rob.scala:310:28
        rob_uop_1_1_pc_lob = _RANDOM[11'h1C3][16:11];	// rob.scala:310:28
        rob_uop_1_1_pdst = _RANDOM[11'h1C5][11:5];	// rob.scala:310:28
        rob_uop_1_1_stale_pdst = _RANDOM[11'h1C6][16:10];	// rob.scala:310:28
        rob_uop_1_1_is_fencei = _RANDOM[11'h1C8][28];	// rob.scala:310:28
        rob_uop_1_1_uses_ldq = _RANDOM[11'h1C8][30];	// rob.scala:310:28
        rob_uop_1_1_uses_stq = _RANDOM[11'h1C8][31];	// rob.scala:310:28
        rob_uop_1_1_is_sys_pc2epc = _RANDOM[11'h1C9][0];	// rob.scala:310:28
        rob_uop_1_1_flush_on_commit = _RANDOM[11'h1C9][2];	// rob.scala:310:28
        rob_uop_1_1_ldst = _RANDOM[11'h1C9][9:4];	// rob.scala:310:28
        rob_uop_1_1_ldst_val = _RANDOM[11'h1C9][28];	// rob.scala:310:28
        rob_uop_1_1_dst_rtype = _RANDOM[11'h1C9][30:29];	// rob.scala:310:28
        rob_uop_1_1_fp_val = _RANDOM[11'h1CA][4];	// rob.scala:310:28
        rob_uop_1_2_uopc = _RANDOM[11'h1CA][21:15];	// rob.scala:310:28
        rob_uop_1_2_is_rvc = _RANDOM[11'h1CC][22];	// rob.scala:310:28
        rob_uop_1_2_br_mask = _RANDOM[11'h1CF][26:11];	// rob.scala:310:28
        rob_uop_1_2_ftq_idx = {_RANDOM[11'h1CF][31], _RANDOM[11'h1D0][3:0]};	// rob.scala:310:28
        rob_uop_1_2_edge_inst = _RANDOM[11'h1D0][4];	// rob.scala:310:28
        rob_uop_1_2_pc_lob = _RANDOM[11'h1D0][10:5];	// rob.scala:310:28
        rob_uop_1_2_pdst = {_RANDOM[11'h1D1][31], _RANDOM[11'h1D2][5:0]};	// rob.scala:310:28
        rob_uop_1_2_stale_pdst = _RANDOM[11'h1D3][10:4];	// rob.scala:310:28
        rob_uop_1_2_is_fencei = _RANDOM[11'h1D5][22];	// rob.scala:310:28
        rob_uop_1_2_uses_ldq = _RANDOM[11'h1D5][24];	// rob.scala:310:28
        rob_uop_1_2_uses_stq = _RANDOM[11'h1D5][25];	// rob.scala:310:28
        rob_uop_1_2_is_sys_pc2epc = _RANDOM[11'h1D5][26];	// rob.scala:310:28
        rob_uop_1_2_flush_on_commit = _RANDOM[11'h1D5][28];	// rob.scala:310:28
        rob_uop_1_2_ldst = {_RANDOM[11'h1D5][31:30], _RANDOM[11'h1D6][3:0]};	// rob.scala:310:28
        rob_uop_1_2_ldst_val = _RANDOM[11'h1D6][22];	// rob.scala:310:28
        rob_uop_1_2_dst_rtype = _RANDOM[11'h1D6][24:23];	// rob.scala:310:28
        rob_uop_1_2_fp_val = _RANDOM[11'h1D6][30];	// rob.scala:310:28
        rob_uop_1_3_uopc = _RANDOM[11'h1D7][15:9];	// rob.scala:310:28
        rob_uop_1_3_is_rvc = _RANDOM[11'h1D9][16];	// rob.scala:310:28
        rob_uop_1_3_br_mask = _RANDOM[11'h1DC][20:5];	// rob.scala:310:28
        rob_uop_1_3_ftq_idx = _RANDOM[11'h1DC][29:25];	// rob.scala:310:28
        rob_uop_1_3_edge_inst = _RANDOM[11'h1DC][30];	// rob.scala:310:28
        rob_uop_1_3_pc_lob = {_RANDOM[11'h1DC][31], _RANDOM[11'h1DD][4:0]};	// rob.scala:310:28
        rob_uop_1_3_pdst = _RANDOM[11'h1DE][31:25];	// rob.scala:310:28
        rob_uop_1_3_stale_pdst = {_RANDOM[11'h1DF][31:30], _RANDOM[11'h1E0][4:0]};	// rob.scala:310:28
        rob_uop_1_3_is_fencei = _RANDOM[11'h1E2][16];	// rob.scala:310:28
        rob_uop_1_3_uses_ldq = _RANDOM[11'h1E2][18];	// rob.scala:310:28
        rob_uop_1_3_uses_stq = _RANDOM[11'h1E2][19];	// rob.scala:310:28
        rob_uop_1_3_is_sys_pc2epc = _RANDOM[11'h1E2][20];	// rob.scala:310:28
        rob_uop_1_3_flush_on_commit = _RANDOM[11'h1E2][22];	// rob.scala:310:28
        rob_uop_1_3_ldst = _RANDOM[11'h1E2][29:24];	// rob.scala:310:28
        rob_uop_1_3_ldst_val = _RANDOM[11'h1E3][16];	// rob.scala:310:28
        rob_uop_1_3_dst_rtype = _RANDOM[11'h1E3][18:17];	// rob.scala:310:28
        rob_uop_1_3_fp_val = _RANDOM[11'h1E3][24];	// rob.scala:310:28
        rob_uop_1_4_uopc = _RANDOM[11'h1E4][9:3];	// rob.scala:310:28
        rob_uop_1_4_is_rvc = _RANDOM[11'h1E6][10];	// rob.scala:310:28
        rob_uop_1_4_br_mask = {_RANDOM[11'h1E8][31], _RANDOM[11'h1E9][14:0]};	// rob.scala:310:28
        rob_uop_1_4_ftq_idx = _RANDOM[11'h1E9][23:19];	// rob.scala:310:28
        rob_uop_1_4_edge_inst = _RANDOM[11'h1E9][24];	// rob.scala:310:28
        rob_uop_1_4_pc_lob = _RANDOM[11'h1E9][30:25];	// rob.scala:310:28
        rob_uop_1_4_pdst = _RANDOM[11'h1EB][25:19];	// rob.scala:310:28
        rob_uop_1_4_stale_pdst = _RANDOM[11'h1EC][30:24];	// rob.scala:310:28
        rob_uop_1_4_is_fencei = _RANDOM[11'h1EF][10];	// rob.scala:310:28
        rob_uop_1_4_uses_ldq = _RANDOM[11'h1EF][12];	// rob.scala:310:28
        rob_uop_1_4_uses_stq = _RANDOM[11'h1EF][13];	// rob.scala:310:28
        rob_uop_1_4_is_sys_pc2epc = _RANDOM[11'h1EF][14];	// rob.scala:310:28
        rob_uop_1_4_flush_on_commit = _RANDOM[11'h1EF][16];	// rob.scala:310:28
        rob_uop_1_4_ldst = _RANDOM[11'h1EF][23:18];	// rob.scala:310:28
        rob_uop_1_4_ldst_val = _RANDOM[11'h1F0][10];	// rob.scala:310:28
        rob_uop_1_4_dst_rtype = _RANDOM[11'h1F0][12:11];	// rob.scala:310:28
        rob_uop_1_4_fp_val = _RANDOM[11'h1F0][18];	// rob.scala:310:28
        rob_uop_1_5_uopc = {_RANDOM[11'h1F0][31:29], _RANDOM[11'h1F1][3:0]};	// rob.scala:310:28
        rob_uop_1_5_is_rvc = _RANDOM[11'h1F3][4];	// rob.scala:310:28
        rob_uop_1_5_br_mask = {_RANDOM[11'h1F5][31:25], _RANDOM[11'h1F6][8:0]};	// rob.scala:310:28
        rob_uop_1_5_ftq_idx = _RANDOM[11'h1F6][17:13];	// rob.scala:310:28
        rob_uop_1_5_edge_inst = _RANDOM[11'h1F6][18];	// rob.scala:310:28
        rob_uop_1_5_pc_lob = _RANDOM[11'h1F6][24:19];	// rob.scala:310:28
        rob_uop_1_5_pdst = _RANDOM[11'h1F8][19:13];	// rob.scala:310:28
        rob_uop_1_5_stale_pdst = _RANDOM[11'h1F9][24:18];	// rob.scala:310:28
        rob_uop_1_5_is_fencei = _RANDOM[11'h1FC][4];	// rob.scala:310:28
        rob_uop_1_5_uses_ldq = _RANDOM[11'h1FC][6];	// rob.scala:310:28
        rob_uop_1_5_uses_stq = _RANDOM[11'h1FC][7];	// rob.scala:310:28
        rob_uop_1_5_is_sys_pc2epc = _RANDOM[11'h1FC][8];	// rob.scala:310:28
        rob_uop_1_5_flush_on_commit = _RANDOM[11'h1FC][10];	// rob.scala:310:28
        rob_uop_1_5_ldst = _RANDOM[11'h1FC][17:12];	// rob.scala:310:28
        rob_uop_1_5_ldst_val = _RANDOM[11'h1FD][4];	// rob.scala:310:28
        rob_uop_1_5_dst_rtype = _RANDOM[11'h1FD][6:5];	// rob.scala:310:28
        rob_uop_1_5_fp_val = _RANDOM[11'h1FD][12];	// rob.scala:310:28
        rob_uop_1_6_uopc = _RANDOM[11'h1FD][29:23];	// rob.scala:310:28
        rob_uop_1_6_is_rvc = _RANDOM[11'h1FF][30];	// rob.scala:310:28
        rob_uop_1_6_br_mask = {_RANDOM[11'h202][31:19], _RANDOM[11'h203][2:0]};	// rob.scala:310:28
        rob_uop_1_6_ftq_idx = _RANDOM[11'h203][11:7];	// rob.scala:310:28
        rob_uop_1_6_edge_inst = _RANDOM[11'h203][12];	// rob.scala:310:28
        rob_uop_1_6_pc_lob = _RANDOM[11'h203][18:13];	// rob.scala:310:28
        rob_uop_1_6_pdst = _RANDOM[11'h205][13:7];	// rob.scala:310:28
        rob_uop_1_6_stale_pdst = _RANDOM[11'h206][18:12];	// rob.scala:310:28
        rob_uop_1_6_is_fencei = _RANDOM[11'h208][30];	// rob.scala:310:28
        rob_uop_1_6_uses_ldq = _RANDOM[11'h209][0];	// rob.scala:310:28
        rob_uop_1_6_uses_stq = _RANDOM[11'h209][1];	// rob.scala:310:28
        rob_uop_1_6_is_sys_pc2epc = _RANDOM[11'h209][2];	// rob.scala:310:28
        rob_uop_1_6_flush_on_commit = _RANDOM[11'h209][4];	// rob.scala:310:28
        rob_uop_1_6_ldst = _RANDOM[11'h209][11:6];	// rob.scala:310:28
        rob_uop_1_6_ldst_val = _RANDOM[11'h209][30];	// rob.scala:310:28
        rob_uop_1_6_dst_rtype = {_RANDOM[11'h209][31], _RANDOM[11'h20A][0]};	// rob.scala:310:28
        rob_uop_1_6_fp_val = _RANDOM[11'h20A][6];	// rob.scala:310:28
        rob_uop_1_7_uopc = _RANDOM[11'h20A][23:17];	// rob.scala:310:28
        rob_uop_1_7_is_rvc = _RANDOM[11'h20C][24];	// rob.scala:310:28
        rob_uop_1_7_br_mask = _RANDOM[11'h20F][28:13];	// rob.scala:310:28
        rob_uop_1_7_ftq_idx = _RANDOM[11'h210][5:1];	// rob.scala:310:28
        rob_uop_1_7_edge_inst = _RANDOM[11'h210][6];	// rob.scala:310:28
        rob_uop_1_7_pc_lob = _RANDOM[11'h210][12:7];	// rob.scala:310:28
        rob_uop_1_7_pdst = _RANDOM[11'h212][7:1];	// rob.scala:310:28
        rob_uop_1_7_stale_pdst = _RANDOM[11'h213][12:6];	// rob.scala:310:28
        rob_uop_1_7_is_fencei = _RANDOM[11'h215][24];	// rob.scala:310:28
        rob_uop_1_7_uses_ldq = _RANDOM[11'h215][26];	// rob.scala:310:28
        rob_uop_1_7_uses_stq = _RANDOM[11'h215][27];	// rob.scala:310:28
        rob_uop_1_7_is_sys_pc2epc = _RANDOM[11'h215][28];	// rob.scala:310:28
        rob_uop_1_7_flush_on_commit = _RANDOM[11'h215][30];	// rob.scala:310:28
        rob_uop_1_7_ldst = _RANDOM[11'h216][5:0];	// rob.scala:310:28
        rob_uop_1_7_ldst_val = _RANDOM[11'h216][24];	// rob.scala:310:28
        rob_uop_1_7_dst_rtype = _RANDOM[11'h216][26:25];	// rob.scala:310:28
        rob_uop_1_7_fp_val = _RANDOM[11'h217][0];	// rob.scala:310:28
        rob_uop_1_8_uopc = _RANDOM[11'h217][17:11];	// rob.scala:310:28
        rob_uop_1_8_is_rvc = _RANDOM[11'h219][18];	// rob.scala:310:28
        rob_uop_1_8_br_mask = _RANDOM[11'h21C][22:7];	// rob.scala:310:28
        rob_uop_1_8_ftq_idx = _RANDOM[11'h21C][31:27];	// rob.scala:310:28
        rob_uop_1_8_edge_inst = _RANDOM[11'h21D][0];	// rob.scala:310:28
        rob_uop_1_8_pc_lob = _RANDOM[11'h21D][6:1];	// rob.scala:310:28
        rob_uop_1_8_pdst = {_RANDOM[11'h21E][31:27], _RANDOM[11'h21F][1:0]};	// rob.scala:310:28
        rob_uop_1_8_stale_pdst = _RANDOM[11'h220][6:0];	// rob.scala:310:28
        rob_uop_1_8_is_fencei = _RANDOM[11'h222][18];	// rob.scala:310:28
        rob_uop_1_8_uses_ldq = _RANDOM[11'h222][20];	// rob.scala:310:28
        rob_uop_1_8_uses_stq = _RANDOM[11'h222][21];	// rob.scala:310:28
        rob_uop_1_8_is_sys_pc2epc = _RANDOM[11'h222][22];	// rob.scala:310:28
        rob_uop_1_8_flush_on_commit = _RANDOM[11'h222][24];	// rob.scala:310:28
        rob_uop_1_8_ldst = _RANDOM[11'h222][31:26];	// rob.scala:310:28
        rob_uop_1_8_ldst_val = _RANDOM[11'h223][18];	// rob.scala:310:28
        rob_uop_1_8_dst_rtype = _RANDOM[11'h223][20:19];	// rob.scala:310:28
        rob_uop_1_8_fp_val = _RANDOM[11'h223][26];	// rob.scala:310:28
        rob_uop_1_9_uopc = _RANDOM[11'h224][11:5];	// rob.scala:310:28
        rob_uop_1_9_is_rvc = _RANDOM[11'h226][12];	// rob.scala:310:28
        rob_uop_1_9_br_mask = _RANDOM[11'h229][16:1];	// rob.scala:310:28
        rob_uop_1_9_ftq_idx = _RANDOM[11'h229][25:21];	// rob.scala:310:28
        rob_uop_1_9_edge_inst = _RANDOM[11'h229][26];	// rob.scala:310:28
        rob_uop_1_9_pc_lob = {_RANDOM[11'h229][31:27], _RANDOM[11'h22A][0]};	// rob.scala:310:28
        rob_uop_1_9_pdst = _RANDOM[11'h22B][27:21];	// rob.scala:310:28
        rob_uop_1_9_stale_pdst = {_RANDOM[11'h22C][31:26], _RANDOM[11'h22D][0]};	// rob.scala:310:28
        rob_uop_1_9_is_fencei = _RANDOM[11'h22F][12];	// rob.scala:310:28
        rob_uop_1_9_uses_ldq = _RANDOM[11'h22F][14];	// rob.scala:310:28
        rob_uop_1_9_uses_stq = _RANDOM[11'h22F][15];	// rob.scala:310:28
        rob_uop_1_9_is_sys_pc2epc = _RANDOM[11'h22F][16];	// rob.scala:310:28
        rob_uop_1_9_flush_on_commit = _RANDOM[11'h22F][18];	// rob.scala:310:28
        rob_uop_1_9_ldst = _RANDOM[11'h22F][25:20];	// rob.scala:310:28
        rob_uop_1_9_ldst_val = _RANDOM[11'h230][12];	// rob.scala:310:28
        rob_uop_1_9_dst_rtype = _RANDOM[11'h230][14:13];	// rob.scala:310:28
        rob_uop_1_9_fp_val = _RANDOM[11'h230][20];	// rob.scala:310:28
        rob_uop_1_10_uopc = {_RANDOM[11'h230][31], _RANDOM[11'h231][5:0]};	// rob.scala:310:28
        rob_uop_1_10_is_rvc = _RANDOM[11'h233][6];	// rob.scala:310:28
        rob_uop_1_10_br_mask = {_RANDOM[11'h235][31:27], _RANDOM[11'h236][10:0]};	// rob.scala:310:28
        rob_uop_1_10_ftq_idx = _RANDOM[11'h236][19:15];	// rob.scala:310:28
        rob_uop_1_10_edge_inst = _RANDOM[11'h236][20];	// rob.scala:310:28
        rob_uop_1_10_pc_lob = _RANDOM[11'h236][26:21];	// rob.scala:310:28
        rob_uop_1_10_pdst = _RANDOM[11'h238][21:15];	// rob.scala:310:28
        rob_uop_1_10_stale_pdst = _RANDOM[11'h239][26:20];	// rob.scala:310:28
        rob_uop_1_10_is_fencei = _RANDOM[11'h23C][6];	// rob.scala:310:28
        rob_uop_1_10_uses_ldq = _RANDOM[11'h23C][8];	// rob.scala:310:28
        rob_uop_1_10_uses_stq = _RANDOM[11'h23C][9];	// rob.scala:310:28
        rob_uop_1_10_is_sys_pc2epc = _RANDOM[11'h23C][10];	// rob.scala:310:28
        rob_uop_1_10_flush_on_commit = _RANDOM[11'h23C][12];	// rob.scala:310:28
        rob_uop_1_10_ldst = _RANDOM[11'h23C][19:14];	// rob.scala:310:28
        rob_uop_1_10_ldst_val = _RANDOM[11'h23D][6];	// rob.scala:310:28
        rob_uop_1_10_dst_rtype = _RANDOM[11'h23D][8:7];	// rob.scala:310:28
        rob_uop_1_10_fp_val = _RANDOM[11'h23D][14];	// rob.scala:310:28
        rob_uop_1_11_uopc = _RANDOM[11'h23D][31:25];	// rob.scala:310:28
        rob_uop_1_11_is_rvc = _RANDOM[11'h240][0];	// rob.scala:310:28
        rob_uop_1_11_br_mask = {_RANDOM[11'h242][31:21], _RANDOM[11'h243][4:0]};	// rob.scala:310:28
        rob_uop_1_11_ftq_idx = _RANDOM[11'h243][13:9];	// rob.scala:310:28
        rob_uop_1_11_edge_inst = _RANDOM[11'h243][14];	// rob.scala:310:28
        rob_uop_1_11_pc_lob = _RANDOM[11'h243][20:15];	// rob.scala:310:28
        rob_uop_1_11_pdst = _RANDOM[11'h245][15:9];	// rob.scala:310:28
        rob_uop_1_11_stale_pdst = _RANDOM[11'h246][20:14];	// rob.scala:310:28
        rob_uop_1_11_is_fencei = _RANDOM[11'h249][0];	// rob.scala:310:28
        rob_uop_1_11_uses_ldq = _RANDOM[11'h249][2];	// rob.scala:310:28
        rob_uop_1_11_uses_stq = _RANDOM[11'h249][3];	// rob.scala:310:28
        rob_uop_1_11_is_sys_pc2epc = _RANDOM[11'h249][4];	// rob.scala:310:28
        rob_uop_1_11_flush_on_commit = _RANDOM[11'h249][6];	// rob.scala:310:28
        rob_uop_1_11_ldst = _RANDOM[11'h249][13:8];	// rob.scala:310:28
        rob_uop_1_11_ldst_val = _RANDOM[11'h24A][0];	// rob.scala:310:28
        rob_uop_1_11_dst_rtype = _RANDOM[11'h24A][2:1];	// rob.scala:310:28
        rob_uop_1_11_fp_val = _RANDOM[11'h24A][8];	// rob.scala:310:28
        rob_uop_1_12_uopc = _RANDOM[11'h24A][25:19];	// rob.scala:310:28
        rob_uop_1_12_is_rvc = _RANDOM[11'h24C][26];	// rob.scala:310:28
        rob_uop_1_12_br_mask = _RANDOM[11'h24F][30:15];	// rob.scala:310:28
        rob_uop_1_12_ftq_idx = _RANDOM[11'h250][7:3];	// rob.scala:310:28
        rob_uop_1_12_edge_inst = _RANDOM[11'h250][8];	// rob.scala:310:28
        rob_uop_1_12_pc_lob = _RANDOM[11'h250][14:9];	// rob.scala:310:28
        rob_uop_1_12_pdst = _RANDOM[11'h252][9:3];	// rob.scala:310:28
        rob_uop_1_12_stale_pdst = _RANDOM[11'h253][14:8];	// rob.scala:310:28
        rob_uop_1_12_is_fencei = _RANDOM[11'h255][26];	// rob.scala:310:28
        rob_uop_1_12_uses_ldq = _RANDOM[11'h255][28];	// rob.scala:310:28
        rob_uop_1_12_uses_stq = _RANDOM[11'h255][29];	// rob.scala:310:28
        rob_uop_1_12_is_sys_pc2epc = _RANDOM[11'h255][30];	// rob.scala:310:28
        rob_uop_1_12_flush_on_commit = _RANDOM[11'h256][0];	// rob.scala:310:28
        rob_uop_1_12_ldst = _RANDOM[11'h256][7:2];	// rob.scala:310:28
        rob_uop_1_12_ldst_val = _RANDOM[11'h256][26];	// rob.scala:310:28
        rob_uop_1_12_dst_rtype = _RANDOM[11'h256][28:27];	// rob.scala:310:28
        rob_uop_1_12_fp_val = _RANDOM[11'h257][2];	// rob.scala:310:28
        rob_uop_1_13_uopc = _RANDOM[11'h257][19:13];	// rob.scala:310:28
        rob_uop_1_13_is_rvc = _RANDOM[11'h259][20];	// rob.scala:310:28
        rob_uop_1_13_br_mask = _RANDOM[11'h25C][24:9];	// rob.scala:310:28
        rob_uop_1_13_ftq_idx = {_RANDOM[11'h25C][31:29], _RANDOM[11'h25D][1:0]};	// rob.scala:310:28
        rob_uop_1_13_edge_inst = _RANDOM[11'h25D][2];	// rob.scala:310:28
        rob_uop_1_13_pc_lob = _RANDOM[11'h25D][8:3];	// rob.scala:310:28
        rob_uop_1_13_pdst = {_RANDOM[11'h25E][31:29], _RANDOM[11'h25F][3:0]};	// rob.scala:310:28
        rob_uop_1_13_stale_pdst = _RANDOM[11'h260][8:2];	// rob.scala:310:28
        rob_uop_1_13_is_fencei = _RANDOM[11'h262][20];	// rob.scala:310:28
        rob_uop_1_13_uses_ldq = _RANDOM[11'h262][22];	// rob.scala:310:28
        rob_uop_1_13_uses_stq = _RANDOM[11'h262][23];	// rob.scala:310:28
        rob_uop_1_13_is_sys_pc2epc = _RANDOM[11'h262][24];	// rob.scala:310:28
        rob_uop_1_13_flush_on_commit = _RANDOM[11'h262][26];	// rob.scala:310:28
        rob_uop_1_13_ldst = {_RANDOM[11'h262][31:28], _RANDOM[11'h263][1:0]};	// rob.scala:310:28
        rob_uop_1_13_ldst_val = _RANDOM[11'h263][20];	// rob.scala:310:28
        rob_uop_1_13_dst_rtype = _RANDOM[11'h263][22:21];	// rob.scala:310:28
        rob_uop_1_13_fp_val = _RANDOM[11'h263][28];	// rob.scala:310:28
        rob_uop_1_14_uopc = _RANDOM[11'h264][13:7];	// rob.scala:310:28
        rob_uop_1_14_is_rvc = _RANDOM[11'h266][14];	// rob.scala:310:28
        rob_uop_1_14_br_mask = _RANDOM[11'h269][18:3];	// rob.scala:310:28
        rob_uop_1_14_ftq_idx = _RANDOM[11'h269][27:23];	// rob.scala:310:28
        rob_uop_1_14_edge_inst = _RANDOM[11'h269][28];	// rob.scala:310:28
        rob_uop_1_14_pc_lob = {_RANDOM[11'h269][31:29], _RANDOM[11'h26A][2:0]};	// rob.scala:310:28
        rob_uop_1_14_pdst = _RANDOM[11'h26B][29:23];	// rob.scala:310:28
        rob_uop_1_14_stale_pdst = {_RANDOM[11'h26C][31:28], _RANDOM[11'h26D][2:0]};	// rob.scala:310:28
        rob_uop_1_14_is_fencei = _RANDOM[11'h26F][14];	// rob.scala:310:28
        rob_uop_1_14_uses_ldq = _RANDOM[11'h26F][16];	// rob.scala:310:28
        rob_uop_1_14_uses_stq = _RANDOM[11'h26F][17];	// rob.scala:310:28
        rob_uop_1_14_is_sys_pc2epc = _RANDOM[11'h26F][18];	// rob.scala:310:28
        rob_uop_1_14_flush_on_commit = _RANDOM[11'h26F][20];	// rob.scala:310:28
        rob_uop_1_14_ldst = _RANDOM[11'h26F][27:22];	// rob.scala:310:28
        rob_uop_1_14_ldst_val = _RANDOM[11'h270][14];	// rob.scala:310:28
        rob_uop_1_14_dst_rtype = _RANDOM[11'h270][16:15];	// rob.scala:310:28
        rob_uop_1_14_fp_val = _RANDOM[11'h270][22];	// rob.scala:310:28
        rob_uop_1_15_uopc = _RANDOM[11'h271][7:1];	// rob.scala:310:28
        rob_uop_1_15_is_rvc = _RANDOM[11'h273][8];	// rob.scala:310:28
        rob_uop_1_15_br_mask = {_RANDOM[11'h275][31:29], _RANDOM[11'h276][12:0]};	// rob.scala:310:28
        rob_uop_1_15_ftq_idx = _RANDOM[11'h276][21:17];	// rob.scala:310:28
        rob_uop_1_15_edge_inst = _RANDOM[11'h276][22];	// rob.scala:310:28
        rob_uop_1_15_pc_lob = _RANDOM[11'h276][28:23];	// rob.scala:310:28
        rob_uop_1_15_pdst = _RANDOM[11'h278][23:17];	// rob.scala:310:28
        rob_uop_1_15_stale_pdst = _RANDOM[11'h279][28:22];	// rob.scala:310:28
        rob_uop_1_15_is_fencei = _RANDOM[11'h27C][8];	// rob.scala:310:28
        rob_uop_1_15_uses_ldq = _RANDOM[11'h27C][10];	// rob.scala:310:28
        rob_uop_1_15_uses_stq = _RANDOM[11'h27C][11];	// rob.scala:310:28
        rob_uop_1_15_is_sys_pc2epc = _RANDOM[11'h27C][12];	// rob.scala:310:28
        rob_uop_1_15_flush_on_commit = _RANDOM[11'h27C][14];	// rob.scala:310:28
        rob_uop_1_15_ldst = _RANDOM[11'h27C][21:16];	// rob.scala:310:28
        rob_uop_1_15_ldst_val = _RANDOM[11'h27D][8];	// rob.scala:310:28
        rob_uop_1_15_dst_rtype = _RANDOM[11'h27D][10:9];	// rob.scala:310:28
        rob_uop_1_15_fp_val = _RANDOM[11'h27D][16];	// rob.scala:310:28
        rob_uop_1_16_uopc = {_RANDOM[11'h27D][31:27], _RANDOM[11'h27E][1:0]};	// rob.scala:310:28
        rob_uop_1_16_is_rvc = _RANDOM[11'h280][2];	// rob.scala:310:28
        rob_uop_1_16_br_mask = {_RANDOM[11'h282][31:23], _RANDOM[11'h283][6:0]};	// rob.scala:310:28
        rob_uop_1_16_ftq_idx = _RANDOM[11'h283][15:11];	// rob.scala:310:28
        rob_uop_1_16_edge_inst = _RANDOM[11'h283][16];	// rob.scala:310:28
        rob_uop_1_16_pc_lob = _RANDOM[11'h283][22:17];	// rob.scala:310:28
        rob_uop_1_16_pdst = _RANDOM[11'h285][17:11];	// rob.scala:310:28
        rob_uop_1_16_stale_pdst = _RANDOM[11'h286][22:16];	// rob.scala:310:28
        rob_uop_1_16_is_fencei = _RANDOM[11'h289][2];	// rob.scala:310:28
        rob_uop_1_16_uses_ldq = _RANDOM[11'h289][4];	// rob.scala:310:28
        rob_uop_1_16_uses_stq = _RANDOM[11'h289][5];	// rob.scala:310:28
        rob_uop_1_16_is_sys_pc2epc = _RANDOM[11'h289][6];	// rob.scala:310:28
        rob_uop_1_16_flush_on_commit = _RANDOM[11'h289][8];	// rob.scala:310:28
        rob_uop_1_16_ldst = _RANDOM[11'h289][15:10];	// rob.scala:310:28
        rob_uop_1_16_ldst_val = _RANDOM[11'h28A][2];	// rob.scala:310:28
        rob_uop_1_16_dst_rtype = _RANDOM[11'h28A][4:3];	// rob.scala:310:28
        rob_uop_1_16_fp_val = _RANDOM[11'h28A][10];	// rob.scala:310:28
        rob_uop_1_17_uopc = _RANDOM[11'h28A][27:21];	// rob.scala:310:28
        rob_uop_1_17_is_rvc = _RANDOM[11'h28C][28];	// rob.scala:310:28
        rob_uop_1_17_br_mask = {_RANDOM[11'h28F][31:17], _RANDOM[11'h290][0]};	// rob.scala:310:28
        rob_uop_1_17_ftq_idx = _RANDOM[11'h290][9:5];	// rob.scala:310:28
        rob_uop_1_17_edge_inst = _RANDOM[11'h290][10];	// rob.scala:310:28
        rob_uop_1_17_pc_lob = _RANDOM[11'h290][16:11];	// rob.scala:310:28
        rob_uop_1_17_pdst = _RANDOM[11'h292][11:5];	// rob.scala:310:28
        rob_uop_1_17_stale_pdst = _RANDOM[11'h293][16:10];	// rob.scala:310:28
        rob_uop_1_17_is_fencei = _RANDOM[11'h295][28];	// rob.scala:310:28
        rob_uop_1_17_uses_ldq = _RANDOM[11'h295][30];	// rob.scala:310:28
        rob_uop_1_17_uses_stq = _RANDOM[11'h295][31];	// rob.scala:310:28
        rob_uop_1_17_is_sys_pc2epc = _RANDOM[11'h296][0];	// rob.scala:310:28
        rob_uop_1_17_flush_on_commit = _RANDOM[11'h296][2];	// rob.scala:310:28
        rob_uop_1_17_ldst = _RANDOM[11'h296][9:4];	// rob.scala:310:28
        rob_uop_1_17_ldst_val = _RANDOM[11'h296][28];	// rob.scala:310:28
        rob_uop_1_17_dst_rtype = _RANDOM[11'h296][30:29];	// rob.scala:310:28
        rob_uop_1_17_fp_val = _RANDOM[11'h297][4];	// rob.scala:310:28
        rob_uop_1_18_uopc = _RANDOM[11'h297][21:15];	// rob.scala:310:28
        rob_uop_1_18_is_rvc = _RANDOM[11'h299][22];	// rob.scala:310:28
        rob_uop_1_18_br_mask = _RANDOM[11'h29C][26:11];	// rob.scala:310:28
        rob_uop_1_18_ftq_idx = {_RANDOM[11'h29C][31], _RANDOM[11'h29D][3:0]};	// rob.scala:310:28
        rob_uop_1_18_edge_inst = _RANDOM[11'h29D][4];	// rob.scala:310:28
        rob_uop_1_18_pc_lob = _RANDOM[11'h29D][10:5];	// rob.scala:310:28
        rob_uop_1_18_pdst = {_RANDOM[11'h29E][31], _RANDOM[11'h29F][5:0]};	// rob.scala:310:28
        rob_uop_1_18_stale_pdst = _RANDOM[11'h2A0][10:4];	// rob.scala:310:28
        rob_uop_1_18_is_fencei = _RANDOM[11'h2A2][22];	// rob.scala:310:28
        rob_uop_1_18_uses_ldq = _RANDOM[11'h2A2][24];	// rob.scala:310:28
        rob_uop_1_18_uses_stq = _RANDOM[11'h2A2][25];	// rob.scala:310:28
        rob_uop_1_18_is_sys_pc2epc = _RANDOM[11'h2A2][26];	// rob.scala:310:28
        rob_uop_1_18_flush_on_commit = _RANDOM[11'h2A2][28];	// rob.scala:310:28
        rob_uop_1_18_ldst = {_RANDOM[11'h2A2][31:30], _RANDOM[11'h2A3][3:0]};	// rob.scala:310:28
        rob_uop_1_18_ldst_val = _RANDOM[11'h2A3][22];	// rob.scala:310:28
        rob_uop_1_18_dst_rtype = _RANDOM[11'h2A3][24:23];	// rob.scala:310:28
        rob_uop_1_18_fp_val = _RANDOM[11'h2A3][30];	// rob.scala:310:28
        rob_uop_1_19_uopc = _RANDOM[11'h2A4][15:9];	// rob.scala:310:28
        rob_uop_1_19_is_rvc = _RANDOM[11'h2A6][16];	// rob.scala:310:28
        rob_uop_1_19_br_mask = _RANDOM[11'h2A9][20:5];	// rob.scala:310:28
        rob_uop_1_19_ftq_idx = _RANDOM[11'h2A9][29:25];	// rob.scala:310:28
        rob_uop_1_19_edge_inst = _RANDOM[11'h2A9][30];	// rob.scala:310:28
        rob_uop_1_19_pc_lob = {_RANDOM[11'h2A9][31], _RANDOM[11'h2AA][4:0]};	// rob.scala:310:28
        rob_uop_1_19_pdst = _RANDOM[11'h2AB][31:25];	// rob.scala:310:28
        rob_uop_1_19_stale_pdst = {_RANDOM[11'h2AC][31:30], _RANDOM[11'h2AD][4:0]};	// rob.scala:310:28
        rob_uop_1_19_is_fencei = _RANDOM[11'h2AF][16];	// rob.scala:310:28
        rob_uop_1_19_uses_ldq = _RANDOM[11'h2AF][18];	// rob.scala:310:28
        rob_uop_1_19_uses_stq = _RANDOM[11'h2AF][19];	// rob.scala:310:28
        rob_uop_1_19_is_sys_pc2epc = _RANDOM[11'h2AF][20];	// rob.scala:310:28
        rob_uop_1_19_flush_on_commit = _RANDOM[11'h2AF][22];	// rob.scala:310:28
        rob_uop_1_19_ldst = _RANDOM[11'h2AF][29:24];	// rob.scala:310:28
        rob_uop_1_19_ldst_val = _RANDOM[11'h2B0][16];	// rob.scala:310:28
        rob_uop_1_19_dst_rtype = _RANDOM[11'h2B0][18:17];	// rob.scala:310:28
        rob_uop_1_19_fp_val = _RANDOM[11'h2B0][24];	// rob.scala:310:28
        rob_uop_1_20_uopc = _RANDOM[11'h2B1][9:3];	// rob.scala:310:28
        rob_uop_1_20_is_rvc = _RANDOM[11'h2B3][10];	// rob.scala:310:28
        rob_uop_1_20_br_mask = {_RANDOM[11'h2B5][31], _RANDOM[11'h2B6][14:0]};	// rob.scala:310:28
        rob_uop_1_20_ftq_idx = _RANDOM[11'h2B6][23:19];	// rob.scala:310:28
        rob_uop_1_20_edge_inst = _RANDOM[11'h2B6][24];	// rob.scala:310:28
        rob_uop_1_20_pc_lob = _RANDOM[11'h2B6][30:25];	// rob.scala:310:28
        rob_uop_1_20_pdst = _RANDOM[11'h2B8][25:19];	// rob.scala:310:28
        rob_uop_1_20_stale_pdst = _RANDOM[11'h2B9][30:24];	// rob.scala:310:28
        rob_uop_1_20_is_fencei = _RANDOM[11'h2BC][10];	// rob.scala:310:28
        rob_uop_1_20_uses_ldq = _RANDOM[11'h2BC][12];	// rob.scala:310:28
        rob_uop_1_20_uses_stq = _RANDOM[11'h2BC][13];	// rob.scala:310:28
        rob_uop_1_20_is_sys_pc2epc = _RANDOM[11'h2BC][14];	// rob.scala:310:28
        rob_uop_1_20_flush_on_commit = _RANDOM[11'h2BC][16];	// rob.scala:310:28
        rob_uop_1_20_ldst = _RANDOM[11'h2BC][23:18];	// rob.scala:310:28
        rob_uop_1_20_ldst_val = _RANDOM[11'h2BD][10];	// rob.scala:310:28
        rob_uop_1_20_dst_rtype = _RANDOM[11'h2BD][12:11];	// rob.scala:310:28
        rob_uop_1_20_fp_val = _RANDOM[11'h2BD][18];	// rob.scala:310:28
        rob_uop_1_21_uopc = {_RANDOM[11'h2BD][31:29], _RANDOM[11'h2BE][3:0]};	// rob.scala:310:28
        rob_uop_1_21_is_rvc = _RANDOM[11'h2C0][4];	// rob.scala:310:28
        rob_uop_1_21_br_mask = {_RANDOM[11'h2C2][31:25], _RANDOM[11'h2C3][8:0]};	// rob.scala:310:28
        rob_uop_1_21_ftq_idx = _RANDOM[11'h2C3][17:13];	// rob.scala:310:28
        rob_uop_1_21_edge_inst = _RANDOM[11'h2C3][18];	// rob.scala:310:28
        rob_uop_1_21_pc_lob = _RANDOM[11'h2C3][24:19];	// rob.scala:310:28
        rob_uop_1_21_pdst = _RANDOM[11'h2C5][19:13];	// rob.scala:310:28
        rob_uop_1_21_stale_pdst = _RANDOM[11'h2C6][24:18];	// rob.scala:310:28
        rob_uop_1_21_is_fencei = _RANDOM[11'h2C9][4];	// rob.scala:310:28
        rob_uop_1_21_uses_ldq = _RANDOM[11'h2C9][6];	// rob.scala:310:28
        rob_uop_1_21_uses_stq = _RANDOM[11'h2C9][7];	// rob.scala:310:28
        rob_uop_1_21_is_sys_pc2epc = _RANDOM[11'h2C9][8];	// rob.scala:310:28
        rob_uop_1_21_flush_on_commit = _RANDOM[11'h2C9][10];	// rob.scala:310:28
        rob_uop_1_21_ldst = _RANDOM[11'h2C9][17:12];	// rob.scala:310:28
        rob_uop_1_21_ldst_val = _RANDOM[11'h2CA][4];	// rob.scala:310:28
        rob_uop_1_21_dst_rtype = _RANDOM[11'h2CA][6:5];	// rob.scala:310:28
        rob_uop_1_21_fp_val = _RANDOM[11'h2CA][12];	// rob.scala:310:28
        rob_uop_1_22_uopc = _RANDOM[11'h2CA][29:23];	// rob.scala:310:28
        rob_uop_1_22_is_rvc = _RANDOM[11'h2CC][30];	// rob.scala:310:28
        rob_uop_1_22_br_mask = {_RANDOM[11'h2CF][31:19], _RANDOM[11'h2D0][2:0]};	// rob.scala:310:28
        rob_uop_1_22_ftq_idx = _RANDOM[11'h2D0][11:7];	// rob.scala:310:28
        rob_uop_1_22_edge_inst = _RANDOM[11'h2D0][12];	// rob.scala:310:28
        rob_uop_1_22_pc_lob = _RANDOM[11'h2D0][18:13];	// rob.scala:310:28
        rob_uop_1_22_pdst = _RANDOM[11'h2D2][13:7];	// rob.scala:310:28
        rob_uop_1_22_stale_pdst = _RANDOM[11'h2D3][18:12];	// rob.scala:310:28
        rob_uop_1_22_is_fencei = _RANDOM[11'h2D5][30];	// rob.scala:310:28
        rob_uop_1_22_uses_ldq = _RANDOM[11'h2D6][0];	// rob.scala:310:28
        rob_uop_1_22_uses_stq = _RANDOM[11'h2D6][1];	// rob.scala:310:28
        rob_uop_1_22_is_sys_pc2epc = _RANDOM[11'h2D6][2];	// rob.scala:310:28
        rob_uop_1_22_flush_on_commit = _RANDOM[11'h2D6][4];	// rob.scala:310:28
        rob_uop_1_22_ldst = _RANDOM[11'h2D6][11:6];	// rob.scala:310:28
        rob_uop_1_22_ldst_val = _RANDOM[11'h2D6][30];	// rob.scala:310:28
        rob_uop_1_22_dst_rtype = {_RANDOM[11'h2D6][31], _RANDOM[11'h2D7][0]};	// rob.scala:310:28
        rob_uop_1_22_fp_val = _RANDOM[11'h2D7][6];	// rob.scala:310:28
        rob_uop_1_23_uopc = _RANDOM[11'h2D7][23:17];	// rob.scala:310:28
        rob_uop_1_23_is_rvc = _RANDOM[11'h2D9][24];	// rob.scala:310:28
        rob_uop_1_23_br_mask = _RANDOM[11'h2DC][28:13];	// rob.scala:310:28
        rob_uop_1_23_ftq_idx = _RANDOM[11'h2DD][5:1];	// rob.scala:310:28
        rob_uop_1_23_edge_inst = _RANDOM[11'h2DD][6];	// rob.scala:310:28
        rob_uop_1_23_pc_lob = _RANDOM[11'h2DD][12:7];	// rob.scala:310:28
        rob_uop_1_23_pdst = _RANDOM[11'h2DF][7:1];	// rob.scala:310:28
        rob_uop_1_23_stale_pdst = _RANDOM[11'h2E0][12:6];	// rob.scala:310:28
        rob_uop_1_23_is_fencei = _RANDOM[11'h2E2][24];	// rob.scala:310:28
        rob_uop_1_23_uses_ldq = _RANDOM[11'h2E2][26];	// rob.scala:310:28
        rob_uop_1_23_uses_stq = _RANDOM[11'h2E2][27];	// rob.scala:310:28
        rob_uop_1_23_is_sys_pc2epc = _RANDOM[11'h2E2][28];	// rob.scala:310:28
        rob_uop_1_23_flush_on_commit = _RANDOM[11'h2E2][30];	// rob.scala:310:28
        rob_uop_1_23_ldst = _RANDOM[11'h2E3][5:0];	// rob.scala:310:28
        rob_uop_1_23_ldst_val = _RANDOM[11'h2E3][24];	// rob.scala:310:28
        rob_uop_1_23_dst_rtype = _RANDOM[11'h2E3][26:25];	// rob.scala:310:28
        rob_uop_1_23_fp_val = _RANDOM[11'h2E4][0];	// rob.scala:310:28
        rob_uop_1_24_uopc = _RANDOM[11'h2E4][17:11];	// rob.scala:310:28
        rob_uop_1_24_is_rvc = _RANDOM[11'h2E6][18];	// rob.scala:310:28
        rob_uop_1_24_br_mask = _RANDOM[11'h2E9][22:7];	// rob.scala:310:28
        rob_uop_1_24_ftq_idx = _RANDOM[11'h2E9][31:27];	// rob.scala:310:28
        rob_uop_1_24_edge_inst = _RANDOM[11'h2EA][0];	// rob.scala:310:28
        rob_uop_1_24_pc_lob = _RANDOM[11'h2EA][6:1];	// rob.scala:310:28
        rob_uop_1_24_pdst = {_RANDOM[11'h2EB][31:27], _RANDOM[11'h2EC][1:0]};	// rob.scala:310:28
        rob_uop_1_24_stale_pdst = _RANDOM[11'h2ED][6:0];	// rob.scala:310:28
        rob_uop_1_24_is_fencei = _RANDOM[11'h2EF][18];	// rob.scala:310:28
        rob_uop_1_24_uses_ldq = _RANDOM[11'h2EF][20];	// rob.scala:310:28
        rob_uop_1_24_uses_stq = _RANDOM[11'h2EF][21];	// rob.scala:310:28
        rob_uop_1_24_is_sys_pc2epc = _RANDOM[11'h2EF][22];	// rob.scala:310:28
        rob_uop_1_24_flush_on_commit = _RANDOM[11'h2EF][24];	// rob.scala:310:28
        rob_uop_1_24_ldst = _RANDOM[11'h2EF][31:26];	// rob.scala:310:28
        rob_uop_1_24_ldst_val = _RANDOM[11'h2F0][18];	// rob.scala:310:28
        rob_uop_1_24_dst_rtype = _RANDOM[11'h2F0][20:19];	// rob.scala:310:28
        rob_uop_1_24_fp_val = _RANDOM[11'h2F0][26];	// rob.scala:310:28
        rob_uop_1_25_uopc = _RANDOM[11'h2F1][11:5];	// rob.scala:310:28
        rob_uop_1_25_is_rvc = _RANDOM[11'h2F3][12];	// rob.scala:310:28
        rob_uop_1_25_br_mask = _RANDOM[11'h2F6][16:1];	// rob.scala:310:28
        rob_uop_1_25_ftq_idx = _RANDOM[11'h2F6][25:21];	// rob.scala:310:28
        rob_uop_1_25_edge_inst = _RANDOM[11'h2F6][26];	// rob.scala:310:28
        rob_uop_1_25_pc_lob = {_RANDOM[11'h2F6][31:27], _RANDOM[11'h2F7][0]};	// rob.scala:310:28
        rob_uop_1_25_pdst = _RANDOM[11'h2F8][27:21];	// rob.scala:310:28
        rob_uop_1_25_stale_pdst = {_RANDOM[11'h2F9][31:26], _RANDOM[11'h2FA][0]};	// rob.scala:310:28
        rob_uop_1_25_is_fencei = _RANDOM[11'h2FC][12];	// rob.scala:310:28
        rob_uop_1_25_uses_ldq = _RANDOM[11'h2FC][14];	// rob.scala:310:28
        rob_uop_1_25_uses_stq = _RANDOM[11'h2FC][15];	// rob.scala:310:28
        rob_uop_1_25_is_sys_pc2epc = _RANDOM[11'h2FC][16];	// rob.scala:310:28
        rob_uop_1_25_flush_on_commit = _RANDOM[11'h2FC][18];	// rob.scala:310:28
        rob_uop_1_25_ldst = _RANDOM[11'h2FC][25:20];	// rob.scala:310:28
        rob_uop_1_25_ldst_val = _RANDOM[11'h2FD][12];	// rob.scala:310:28
        rob_uop_1_25_dst_rtype = _RANDOM[11'h2FD][14:13];	// rob.scala:310:28
        rob_uop_1_25_fp_val = _RANDOM[11'h2FD][20];	// rob.scala:310:28
        rob_uop_1_26_uopc = {_RANDOM[11'h2FD][31], _RANDOM[11'h2FE][5:0]};	// rob.scala:310:28
        rob_uop_1_26_is_rvc = _RANDOM[11'h300][6];	// rob.scala:310:28
        rob_uop_1_26_br_mask = {_RANDOM[11'h302][31:27], _RANDOM[11'h303][10:0]};	// rob.scala:310:28
        rob_uop_1_26_ftq_idx = _RANDOM[11'h303][19:15];	// rob.scala:310:28
        rob_uop_1_26_edge_inst = _RANDOM[11'h303][20];	// rob.scala:310:28
        rob_uop_1_26_pc_lob = _RANDOM[11'h303][26:21];	// rob.scala:310:28
        rob_uop_1_26_pdst = _RANDOM[11'h305][21:15];	// rob.scala:310:28
        rob_uop_1_26_stale_pdst = _RANDOM[11'h306][26:20];	// rob.scala:310:28
        rob_uop_1_26_is_fencei = _RANDOM[11'h309][6];	// rob.scala:310:28
        rob_uop_1_26_uses_ldq = _RANDOM[11'h309][8];	// rob.scala:310:28
        rob_uop_1_26_uses_stq = _RANDOM[11'h309][9];	// rob.scala:310:28
        rob_uop_1_26_is_sys_pc2epc = _RANDOM[11'h309][10];	// rob.scala:310:28
        rob_uop_1_26_flush_on_commit = _RANDOM[11'h309][12];	// rob.scala:310:28
        rob_uop_1_26_ldst = _RANDOM[11'h309][19:14];	// rob.scala:310:28
        rob_uop_1_26_ldst_val = _RANDOM[11'h30A][6];	// rob.scala:310:28
        rob_uop_1_26_dst_rtype = _RANDOM[11'h30A][8:7];	// rob.scala:310:28
        rob_uop_1_26_fp_val = _RANDOM[11'h30A][14];	// rob.scala:310:28
        rob_uop_1_27_uopc = _RANDOM[11'h30A][31:25];	// rob.scala:310:28
        rob_uop_1_27_is_rvc = _RANDOM[11'h30D][0];	// rob.scala:310:28
        rob_uop_1_27_br_mask = {_RANDOM[11'h30F][31:21], _RANDOM[11'h310][4:0]};	// rob.scala:310:28
        rob_uop_1_27_ftq_idx = _RANDOM[11'h310][13:9];	// rob.scala:310:28
        rob_uop_1_27_edge_inst = _RANDOM[11'h310][14];	// rob.scala:310:28
        rob_uop_1_27_pc_lob = _RANDOM[11'h310][20:15];	// rob.scala:310:28
        rob_uop_1_27_pdst = _RANDOM[11'h312][15:9];	// rob.scala:310:28
        rob_uop_1_27_stale_pdst = _RANDOM[11'h313][20:14];	// rob.scala:310:28
        rob_uop_1_27_is_fencei = _RANDOM[11'h316][0];	// rob.scala:310:28
        rob_uop_1_27_uses_ldq = _RANDOM[11'h316][2];	// rob.scala:310:28
        rob_uop_1_27_uses_stq = _RANDOM[11'h316][3];	// rob.scala:310:28
        rob_uop_1_27_is_sys_pc2epc = _RANDOM[11'h316][4];	// rob.scala:310:28
        rob_uop_1_27_flush_on_commit = _RANDOM[11'h316][6];	// rob.scala:310:28
        rob_uop_1_27_ldst = _RANDOM[11'h316][13:8];	// rob.scala:310:28
        rob_uop_1_27_ldst_val = _RANDOM[11'h317][0];	// rob.scala:310:28
        rob_uop_1_27_dst_rtype = _RANDOM[11'h317][2:1];	// rob.scala:310:28
        rob_uop_1_27_fp_val = _RANDOM[11'h317][8];	// rob.scala:310:28
        rob_uop_1_28_uopc = _RANDOM[11'h317][25:19];	// rob.scala:310:28
        rob_uop_1_28_is_rvc = _RANDOM[11'h319][26];	// rob.scala:310:28
        rob_uop_1_28_br_mask = _RANDOM[11'h31C][30:15];	// rob.scala:310:28
        rob_uop_1_28_ftq_idx = _RANDOM[11'h31D][7:3];	// rob.scala:310:28
        rob_uop_1_28_edge_inst = _RANDOM[11'h31D][8];	// rob.scala:310:28
        rob_uop_1_28_pc_lob = _RANDOM[11'h31D][14:9];	// rob.scala:310:28
        rob_uop_1_28_pdst = _RANDOM[11'h31F][9:3];	// rob.scala:310:28
        rob_uop_1_28_stale_pdst = _RANDOM[11'h320][14:8];	// rob.scala:310:28
        rob_uop_1_28_is_fencei = _RANDOM[11'h322][26];	// rob.scala:310:28
        rob_uop_1_28_uses_ldq = _RANDOM[11'h322][28];	// rob.scala:310:28
        rob_uop_1_28_uses_stq = _RANDOM[11'h322][29];	// rob.scala:310:28
        rob_uop_1_28_is_sys_pc2epc = _RANDOM[11'h322][30];	// rob.scala:310:28
        rob_uop_1_28_flush_on_commit = _RANDOM[11'h323][0];	// rob.scala:310:28
        rob_uop_1_28_ldst = _RANDOM[11'h323][7:2];	// rob.scala:310:28
        rob_uop_1_28_ldst_val = _RANDOM[11'h323][26];	// rob.scala:310:28
        rob_uop_1_28_dst_rtype = _RANDOM[11'h323][28:27];	// rob.scala:310:28
        rob_uop_1_28_fp_val = _RANDOM[11'h324][2];	// rob.scala:310:28
        rob_uop_1_29_uopc = _RANDOM[11'h324][19:13];	// rob.scala:310:28
        rob_uop_1_29_is_rvc = _RANDOM[11'h326][20];	// rob.scala:310:28
        rob_uop_1_29_br_mask = _RANDOM[11'h329][24:9];	// rob.scala:310:28
        rob_uop_1_29_ftq_idx = {_RANDOM[11'h329][31:29], _RANDOM[11'h32A][1:0]};	// rob.scala:310:28
        rob_uop_1_29_edge_inst = _RANDOM[11'h32A][2];	// rob.scala:310:28
        rob_uop_1_29_pc_lob = _RANDOM[11'h32A][8:3];	// rob.scala:310:28
        rob_uop_1_29_pdst = {_RANDOM[11'h32B][31:29], _RANDOM[11'h32C][3:0]};	// rob.scala:310:28
        rob_uop_1_29_stale_pdst = _RANDOM[11'h32D][8:2];	// rob.scala:310:28
        rob_uop_1_29_is_fencei = _RANDOM[11'h32F][20];	// rob.scala:310:28
        rob_uop_1_29_uses_ldq = _RANDOM[11'h32F][22];	// rob.scala:310:28
        rob_uop_1_29_uses_stq = _RANDOM[11'h32F][23];	// rob.scala:310:28
        rob_uop_1_29_is_sys_pc2epc = _RANDOM[11'h32F][24];	// rob.scala:310:28
        rob_uop_1_29_flush_on_commit = _RANDOM[11'h32F][26];	// rob.scala:310:28
        rob_uop_1_29_ldst = {_RANDOM[11'h32F][31:28], _RANDOM[11'h330][1:0]};	// rob.scala:310:28
        rob_uop_1_29_ldst_val = _RANDOM[11'h330][20];	// rob.scala:310:28
        rob_uop_1_29_dst_rtype = _RANDOM[11'h330][22:21];	// rob.scala:310:28
        rob_uop_1_29_fp_val = _RANDOM[11'h330][28];	// rob.scala:310:28
        rob_uop_1_30_uopc = _RANDOM[11'h331][13:7];	// rob.scala:310:28
        rob_uop_1_30_is_rvc = _RANDOM[11'h333][14];	// rob.scala:310:28
        rob_uop_1_30_br_mask = _RANDOM[11'h336][18:3];	// rob.scala:310:28
        rob_uop_1_30_ftq_idx = _RANDOM[11'h336][27:23];	// rob.scala:310:28
        rob_uop_1_30_edge_inst = _RANDOM[11'h336][28];	// rob.scala:310:28
        rob_uop_1_30_pc_lob = {_RANDOM[11'h336][31:29], _RANDOM[11'h337][2:0]};	// rob.scala:310:28
        rob_uop_1_30_pdst = _RANDOM[11'h338][29:23];	// rob.scala:310:28
        rob_uop_1_30_stale_pdst = {_RANDOM[11'h339][31:28], _RANDOM[11'h33A][2:0]};	// rob.scala:310:28
        rob_uop_1_30_is_fencei = _RANDOM[11'h33C][14];	// rob.scala:310:28
        rob_uop_1_30_uses_ldq = _RANDOM[11'h33C][16];	// rob.scala:310:28
        rob_uop_1_30_uses_stq = _RANDOM[11'h33C][17];	// rob.scala:310:28
        rob_uop_1_30_is_sys_pc2epc = _RANDOM[11'h33C][18];	// rob.scala:310:28
        rob_uop_1_30_flush_on_commit = _RANDOM[11'h33C][20];	// rob.scala:310:28
        rob_uop_1_30_ldst = _RANDOM[11'h33C][27:22];	// rob.scala:310:28
        rob_uop_1_30_ldst_val = _RANDOM[11'h33D][14];	// rob.scala:310:28
        rob_uop_1_30_dst_rtype = _RANDOM[11'h33D][16:15];	// rob.scala:310:28
        rob_uop_1_30_fp_val = _RANDOM[11'h33D][22];	// rob.scala:310:28
        rob_uop_1_31_uopc = _RANDOM[11'h33E][7:1];	// rob.scala:310:28
        rob_uop_1_31_is_rvc = _RANDOM[11'h340][8];	// rob.scala:310:28
        rob_uop_1_31_br_mask = {_RANDOM[11'h342][31:29], _RANDOM[11'h343][12:0]};	// rob.scala:310:28
        rob_uop_1_31_ftq_idx = _RANDOM[11'h343][21:17];	// rob.scala:310:28
        rob_uop_1_31_edge_inst = _RANDOM[11'h343][22];	// rob.scala:310:28
        rob_uop_1_31_pc_lob = _RANDOM[11'h343][28:23];	// rob.scala:310:28
        rob_uop_1_31_pdst = _RANDOM[11'h345][23:17];	// rob.scala:310:28
        rob_uop_1_31_stale_pdst = _RANDOM[11'h346][28:22];	// rob.scala:310:28
        rob_uop_1_31_is_fencei = _RANDOM[11'h349][8];	// rob.scala:310:28
        rob_uop_1_31_uses_ldq = _RANDOM[11'h349][10];	// rob.scala:310:28
        rob_uop_1_31_uses_stq = _RANDOM[11'h349][11];	// rob.scala:310:28
        rob_uop_1_31_is_sys_pc2epc = _RANDOM[11'h349][12];	// rob.scala:310:28
        rob_uop_1_31_flush_on_commit = _RANDOM[11'h349][14];	// rob.scala:310:28
        rob_uop_1_31_ldst = _RANDOM[11'h349][21:16];	// rob.scala:310:28
        rob_uop_1_31_ldst_val = _RANDOM[11'h34A][8];	// rob.scala:310:28
        rob_uop_1_31_dst_rtype = _RANDOM[11'h34A][10:9];	// rob.scala:310:28
        rob_uop_1_31_fp_val = _RANDOM[11'h34A][16];	// rob.scala:310:28
        rob_exception_1_0 = _RANDOM[11'h34A][27];	// rob.scala:310:28, :311:28
        rob_exception_1_1 = _RANDOM[11'h34A][28];	// rob.scala:310:28, :311:28
        rob_exception_1_2 = _RANDOM[11'h34A][29];	// rob.scala:310:28, :311:28
        rob_exception_1_3 = _RANDOM[11'h34A][30];	// rob.scala:310:28, :311:28
        rob_exception_1_4 = _RANDOM[11'h34A][31];	// rob.scala:310:28, :311:28
        rob_exception_1_5 = _RANDOM[11'h34B][0];	// rob.scala:311:28
        rob_exception_1_6 = _RANDOM[11'h34B][1];	// rob.scala:311:28
        rob_exception_1_7 = _RANDOM[11'h34B][2];	// rob.scala:311:28
        rob_exception_1_8 = _RANDOM[11'h34B][3];	// rob.scala:311:28
        rob_exception_1_9 = _RANDOM[11'h34B][4];	// rob.scala:311:28
        rob_exception_1_10 = _RANDOM[11'h34B][5];	// rob.scala:311:28
        rob_exception_1_11 = _RANDOM[11'h34B][6];	// rob.scala:311:28
        rob_exception_1_12 = _RANDOM[11'h34B][7];	// rob.scala:311:28
        rob_exception_1_13 = _RANDOM[11'h34B][8];	// rob.scala:311:28
        rob_exception_1_14 = _RANDOM[11'h34B][9];	// rob.scala:311:28
        rob_exception_1_15 = _RANDOM[11'h34B][10];	// rob.scala:311:28
        rob_exception_1_16 = _RANDOM[11'h34B][11];	// rob.scala:311:28
        rob_exception_1_17 = _RANDOM[11'h34B][12];	// rob.scala:311:28
        rob_exception_1_18 = _RANDOM[11'h34B][13];	// rob.scala:311:28
        rob_exception_1_19 = _RANDOM[11'h34B][14];	// rob.scala:311:28
        rob_exception_1_20 = _RANDOM[11'h34B][15];	// rob.scala:311:28
        rob_exception_1_21 = _RANDOM[11'h34B][16];	// rob.scala:311:28
        rob_exception_1_22 = _RANDOM[11'h34B][17];	// rob.scala:311:28
        rob_exception_1_23 = _RANDOM[11'h34B][18];	// rob.scala:311:28
        rob_exception_1_24 = _RANDOM[11'h34B][19];	// rob.scala:311:28
        rob_exception_1_25 = _RANDOM[11'h34B][20];	// rob.scala:311:28
        rob_exception_1_26 = _RANDOM[11'h34B][21];	// rob.scala:311:28
        rob_exception_1_27 = _RANDOM[11'h34B][22];	// rob.scala:311:28
        rob_exception_1_28 = _RANDOM[11'h34B][23];	// rob.scala:311:28
        rob_exception_1_29 = _RANDOM[11'h34B][24];	// rob.scala:311:28
        rob_exception_1_30 = _RANDOM[11'h34B][25];	// rob.scala:311:28
        rob_exception_1_31 = _RANDOM[11'h34B][26];	// rob.scala:311:28
        rob_predicated_1_0 = _RANDOM[11'h34B][27];	// rob.scala:311:28, :312:29
        rob_predicated_1_1 = _RANDOM[11'h34B][28];	// rob.scala:311:28, :312:29
        rob_predicated_1_2 = _RANDOM[11'h34B][29];	// rob.scala:311:28, :312:29
        rob_predicated_1_3 = _RANDOM[11'h34B][30];	// rob.scala:311:28, :312:29
        rob_predicated_1_4 = _RANDOM[11'h34B][31];	// rob.scala:311:28, :312:29
        rob_predicated_1_5 = _RANDOM[11'h34C][0];	// rob.scala:312:29
        rob_predicated_1_6 = _RANDOM[11'h34C][1];	// rob.scala:312:29
        rob_predicated_1_7 = _RANDOM[11'h34C][2];	// rob.scala:312:29
        rob_predicated_1_8 = _RANDOM[11'h34C][3];	// rob.scala:312:29
        rob_predicated_1_9 = _RANDOM[11'h34C][4];	// rob.scala:312:29
        rob_predicated_1_10 = _RANDOM[11'h34C][5];	// rob.scala:312:29
        rob_predicated_1_11 = _RANDOM[11'h34C][6];	// rob.scala:312:29
        rob_predicated_1_12 = _RANDOM[11'h34C][7];	// rob.scala:312:29
        rob_predicated_1_13 = _RANDOM[11'h34C][8];	// rob.scala:312:29
        rob_predicated_1_14 = _RANDOM[11'h34C][9];	// rob.scala:312:29
        rob_predicated_1_15 = _RANDOM[11'h34C][10];	// rob.scala:312:29
        rob_predicated_1_16 = _RANDOM[11'h34C][11];	// rob.scala:312:29
        rob_predicated_1_17 = _RANDOM[11'h34C][12];	// rob.scala:312:29
        rob_predicated_1_18 = _RANDOM[11'h34C][13];	// rob.scala:312:29
        rob_predicated_1_19 = _RANDOM[11'h34C][14];	// rob.scala:312:29
        rob_predicated_1_20 = _RANDOM[11'h34C][15];	// rob.scala:312:29
        rob_predicated_1_21 = _RANDOM[11'h34C][16];	// rob.scala:312:29
        rob_predicated_1_22 = _RANDOM[11'h34C][17];	// rob.scala:312:29
        rob_predicated_1_23 = _RANDOM[11'h34C][18];	// rob.scala:312:29
        rob_predicated_1_24 = _RANDOM[11'h34C][19];	// rob.scala:312:29
        rob_predicated_1_25 = _RANDOM[11'h34C][20];	// rob.scala:312:29
        rob_predicated_1_26 = _RANDOM[11'h34C][21];	// rob.scala:312:29
        rob_predicated_1_27 = _RANDOM[11'h34C][22];	// rob.scala:312:29
        rob_predicated_1_28 = _RANDOM[11'h34C][23];	// rob.scala:312:29
        rob_predicated_1_29 = _RANDOM[11'h34C][24];	// rob.scala:312:29
        rob_predicated_1_30 = _RANDOM[11'h34C][25];	// rob.scala:312:29
        rob_predicated_1_31 = _RANDOM[11'h34C][26];	// rob.scala:312:29
        rob_val_2_0 = _RANDOM[11'h34C][27];	// rob.scala:307:32, :312:29
        rob_val_2_1 = _RANDOM[11'h34C][28];	// rob.scala:307:32, :312:29
        rob_val_2_2 = _RANDOM[11'h34C][29];	// rob.scala:307:32, :312:29
        rob_val_2_3 = _RANDOM[11'h34C][30];	// rob.scala:307:32, :312:29
        rob_val_2_4 = _RANDOM[11'h34C][31];	// rob.scala:307:32, :312:29
        rob_val_2_5 = _RANDOM[11'h34D][0];	// rob.scala:307:32
        rob_val_2_6 = _RANDOM[11'h34D][1];	// rob.scala:307:32
        rob_val_2_7 = _RANDOM[11'h34D][2];	// rob.scala:307:32
        rob_val_2_8 = _RANDOM[11'h34D][3];	// rob.scala:307:32
        rob_val_2_9 = _RANDOM[11'h34D][4];	// rob.scala:307:32
        rob_val_2_10 = _RANDOM[11'h34D][5];	// rob.scala:307:32
        rob_val_2_11 = _RANDOM[11'h34D][6];	// rob.scala:307:32
        rob_val_2_12 = _RANDOM[11'h34D][7];	// rob.scala:307:32
        rob_val_2_13 = _RANDOM[11'h34D][8];	// rob.scala:307:32
        rob_val_2_14 = _RANDOM[11'h34D][9];	// rob.scala:307:32
        rob_val_2_15 = _RANDOM[11'h34D][10];	// rob.scala:307:32
        rob_val_2_16 = _RANDOM[11'h34D][11];	// rob.scala:307:32
        rob_val_2_17 = _RANDOM[11'h34D][12];	// rob.scala:307:32
        rob_val_2_18 = _RANDOM[11'h34D][13];	// rob.scala:307:32
        rob_val_2_19 = _RANDOM[11'h34D][14];	// rob.scala:307:32
        rob_val_2_20 = _RANDOM[11'h34D][15];	// rob.scala:307:32
        rob_val_2_21 = _RANDOM[11'h34D][16];	// rob.scala:307:32
        rob_val_2_22 = _RANDOM[11'h34D][17];	// rob.scala:307:32
        rob_val_2_23 = _RANDOM[11'h34D][18];	// rob.scala:307:32
        rob_val_2_24 = _RANDOM[11'h34D][19];	// rob.scala:307:32
        rob_val_2_25 = _RANDOM[11'h34D][20];	// rob.scala:307:32
        rob_val_2_26 = _RANDOM[11'h34D][21];	// rob.scala:307:32
        rob_val_2_27 = _RANDOM[11'h34D][22];	// rob.scala:307:32
        rob_val_2_28 = _RANDOM[11'h34D][23];	// rob.scala:307:32
        rob_val_2_29 = _RANDOM[11'h34D][24];	// rob.scala:307:32
        rob_val_2_30 = _RANDOM[11'h34D][25];	// rob.scala:307:32
        rob_val_2_31 = _RANDOM[11'h34D][26];	// rob.scala:307:32
        rob_bsy_2_0 = _RANDOM[11'h34D][27];	// rob.scala:307:32, :308:28
        rob_bsy_2_1 = _RANDOM[11'h34D][28];	// rob.scala:307:32, :308:28
        rob_bsy_2_2 = _RANDOM[11'h34D][29];	// rob.scala:307:32, :308:28
        rob_bsy_2_3 = _RANDOM[11'h34D][30];	// rob.scala:307:32, :308:28
        rob_bsy_2_4 = _RANDOM[11'h34D][31];	// rob.scala:307:32, :308:28
        rob_bsy_2_5 = _RANDOM[11'h34E][0];	// rob.scala:308:28
        rob_bsy_2_6 = _RANDOM[11'h34E][1];	// rob.scala:308:28
        rob_bsy_2_7 = _RANDOM[11'h34E][2];	// rob.scala:308:28
        rob_bsy_2_8 = _RANDOM[11'h34E][3];	// rob.scala:308:28
        rob_bsy_2_9 = _RANDOM[11'h34E][4];	// rob.scala:308:28
        rob_bsy_2_10 = _RANDOM[11'h34E][5];	// rob.scala:308:28
        rob_bsy_2_11 = _RANDOM[11'h34E][6];	// rob.scala:308:28
        rob_bsy_2_12 = _RANDOM[11'h34E][7];	// rob.scala:308:28
        rob_bsy_2_13 = _RANDOM[11'h34E][8];	// rob.scala:308:28
        rob_bsy_2_14 = _RANDOM[11'h34E][9];	// rob.scala:308:28
        rob_bsy_2_15 = _RANDOM[11'h34E][10];	// rob.scala:308:28
        rob_bsy_2_16 = _RANDOM[11'h34E][11];	// rob.scala:308:28
        rob_bsy_2_17 = _RANDOM[11'h34E][12];	// rob.scala:308:28
        rob_bsy_2_18 = _RANDOM[11'h34E][13];	// rob.scala:308:28
        rob_bsy_2_19 = _RANDOM[11'h34E][14];	// rob.scala:308:28
        rob_bsy_2_20 = _RANDOM[11'h34E][15];	// rob.scala:308:28
        rob_bsy_2_21 = _RANDOM[11'h34E][16];	// rob.scala:308:28
        rob_bsy_2_22 = _RANDOM[11'h34E][17];	// rob.scala:308:28
        rob_bsy_2_23 = _RANDOM[11'h34E][18];	// rob.scala:308:28
        rob_bsy_2_24 = _RANDOM[11'h34E][19];	// rob.scala:308:28
        rob_bsy_2_25 = _RANDOM[11'h34E][20];	// rob.scala:308:28
        rob_bsy_2_26 = _RANDOM[11'h34E][21];	// rob.scala:308:28
        rob_bsy_2_27 = _RANDOM[11'h34E][22];	// rob.scala:308:28
        rob_bsy_2_28 = _RANDOM[11'h34E][23];	// rob.scala:308:28
        rob_bsy_2_29 = _RANDOM[11'h34E][24];	// rob.scala:308:28
        rob_bsy_2_30 = _RANDOM[11'h34E][25];	// rob.scala:308:28
        rob_bsy_2_31 = _RANDOM[11'h34E][26];	// rob.scala:308:28
        rob_unsafe_2_0 = _RANDOM[11'h34E][27];	// rob.scala:308:28, :309:28
        rob_unsafe_2_1 = _RANDOM[11'h34E][28];	// rob.scala:308:28, :309:28
        rob_unsafe_2_2 = _RANDOM[11'h34E][29];	// rob.scala:308:28, :309:28
        rob_unsafe_2_3 = _RANDOM[11'h34E][30];	// rob.scala:308:28, :309:28
        rob_unsafe_2_4 = _RANDOM[11'h34E][31];	// rob.scala:308:28, :309:28
        rob_unsafe_2_5 = _RANDOM[11'h34F][0];	// rob.scala:309:28
        rob_unsafe_2_6 = _RANDOM[11'h34F][1];	// rob.scala:309:28
        rob_unsafe_2_7 = _RANDOM[11'h34F][2];	// rob.scala:309:28
        rob_unsafe_2_8 = _RANDOM[11'h34F][3];	// rob.scala:309:28
        rob_unsafe_2_9 = _RANDOM[11'h34F][4];	// rob.scala:309:28
        rob_unsafe_2_10 = _RANDOM[11'h34F][5];	// rob.scala:309:28
        rob_unsafe_2_11 = _RANDOM[11'h34F][6];	// rob.scala:309:28
        rob_unsafe_2_12 = _RANDOM[11'h34F][7];	// rob.scala:309:28
        rob_unsafe_2_13 = _RANDOM[11'h34F][8];	// rob.scala:309:28
        rob_unsafe_2_14 = _RANDOM[11'h34F][9];	// rob.scala:309:28
        rob_unsafe_2_15 = _RANDOM[11'h34F][10];	// rob.scala:309:28
        rob_unsafe_2_16 = _RANDOM[11'h34F][11];	// rob.scala:309:28
        rob_unsafe_2_17 = _RANDOM[11'h34F][12];	// rob.scala:309:28
        rob_unsafe_2_18 = _RANDOM[11'h34F][13];	// rob.scala:309:28
        rob_unsafe_2_19 = _RANDOM[11'h34F][14];	// rob.scala:309:28
        rob_unsafe_2_20 = _RANDOM[11'h34F][15];	// rob.scala:309:28
        rob_unsafe_2_21 = _RANDOM[11'h34F][16];	// rob.scala:309:28
        rob_unsafe_2_22 = _RANDOM[11'h34F][17];	// rob.scala:309:28
        rob_unsafe_2_23 = _RANDOM[11'h34F][18];	// rob.scala:309:28
        rob_unsafe_2_24 = _RANDOM[11'h34F][19];	// rob.scala:309:28
        rob_unsafe_2_25 = _RANDOM[11'h34F][20];	// rob.scala:309:28
        rob_unsafe_2_26 = _RANDOM[11'h34F][21];	// rob.scala:309:28
        rob_unsafe_2_27 = _RANDOM[11'h34F][22];	// rob.scala:309:28
        rob_unsafe_2_28 = _RANDOM[11'h34F][23];	// rob.scala:309:28
        rob_unsafe_2_29 = _RANDOM[11'h34F][24];	// rob.scala:309:28
        rob_unsafe_2_30 = _RANDOM[11'h34F][25];	// rob.scala:309:28
        rob_unsafe_2_31 = _RANDOM[11'h34F][26];	// rob.scala:309:28
        rob_uop_2_0_uopc = {_RANDOM[11'h34F][31:27], _RANDOM[11'h350][1:0]};	// rob.scala:309:28, :310:28
        rob_uop_2_0_is_rvc = _RANDOM[11'h352][2];	// rob.scala:310:28
        rob_uop_2_0_br_mask = {_RANDOM[11'h354][31:23], _RANDOM[11'h355][6:0]};	// rob.scala:310:28
        rob_uop_2_0_ftq_idx = _RANDOM[11'h355][15:11];	// rob.scala:310:28
        rob_uop_2_0_edge_inst = _RANDOM[11'h355][16];	// rob.scala:310:28
        rob_uop_2_0_pc_lob = _RANDOM[11'h355][22:17];	// rob.scala:310:28
        rob_uop_2_0_pdst = _RANDOM[11'h357][17:11];	// rob.scala:310:28
        rob_uop_2_0_stale_pdst = _RANDOM[11'h358][22:16];	// rob.scala:310:28
        rob_uop_2_0_is_fencei = _RANDOM[11'h35B][2];	// rob.scala:310:28
        rob_uop_2_0_uses_ldq = _RANDOM[11'h35B][4];	// rob.scala:310:28
        rob_uop_2_0_uses_stq = _RANDOM[11'h35B][5];	// rob.scala:310:28
        rob_uop_2_0_is_sys_pc2epc = _RANDOM[11'h35B][6];	// rob.scala:310:28
        rob_uop_2_0_flush_on_commit = _RANDOM[11'h35B][8];	// rob.scala:310:28
        rob_uop_2_0_ldst = _RANDOM[11'h35B][15:10];	// rob.scala:310:28
        rob_uop_2_0_ldst_val = _RANDOM[11'h35C][2];	// rob.scala:310:28
        rob_uop_2_0_dst_rtype = _RANDOM[11'h35C][4:3];	// rob.scala:310:28
        rob_uop_2_0_fp_val = _RANDOM[11'h35C][10];	// rob.scala:310:28
        rob_uop_2_1_uopc = _RANDOM[11'h35C][27:21];	// rob.scala:310:28
        rob_uop_2_1_is_rvc = _RANDOM[11'h35E][28];	// rob.scala:310:28
        rob_uop_2_1_br_mask = {_RANDOM[11'h361][31:17], _RANDOM[11'h362][0]};	// rob.scala:310:28
        rob_uop_2_1_ftq_idx = _RANDOM[11'h362][9:5];	// rob.scala:310:28
        rob_uop_2_1_edge_inst = _RANDOM[11'h362][10];	// rob.scala:310:28
        rob_uop_2_1_pc_lob = _RANDOM[11'h362][16:11];	// rob.scala:310:28
        rob_uop_2_1_pdst = _RANDOM[11'h364][11:5];	// rob.scala:310:28
        rob_uop_2_1_stale_pdst = _RANDOM[11'h365][16:10];	// rob.scala:310:28
        rob_uop_2_1_is_fencei = _RANDOM[11'h367][28];	// rob.scala:310:28
        rob_uop_2_1_uses_ldq = _RANDOM[11'h367][30];	// rob.scala:310:28
        rob_uop_2_1_uses_stq = _RANDOM[11'h367][31];	// rob.scala:310:28
        rob_uop_2_1_is_sys_pc2epc = _RANDOM[11'h368][0];	// rob.scala:310:28
        rob_uop_2_1_flush_on_commit = _RANDOM[11'h368][2];	// rob.scala:310:28
        rob_uop_2_1_ldst = _RANDOM[11'h368][9:4];	// rob.scala:310:28
        rob_uop_2_1_ldst_val = _RANDOM[11'h368][28];	// rob.scala:310:28
        rob_uop_2_1_dst_rtype = _RANDOM[11'h368][30:29];	// rob.scala:310:28
        rob_uop_2_1_fp_val = _RANDOM[11'h369][4];	// rob.scala:310:28
        rob_uop_2_2_uopc = _RANDOM[11'h369][21:15];	// rob.scala:310:28
        rob_uop_2_2_is_rvc = _RANDOM[11'h36B][22];	// rob.scala:310:28
        rob_uop_2_2_br_mask = _RANDOM[11'h36E][26:11];	// rob.scala:310:28
        rob_uop_2_2_ftq_idx = {_RANDOM[11'h36E][31], _RANDOM[11'h36F][3:0]};	// rob.scala:310:28
        rob_uop_2_2_edge_inst = _RANDOM[11'h36F][4];	// rob.scala:310:28
        rob_uop_2_2_pc_lob = _RANDOM[11'h36F][10:5];	// rob.scala:310:28
        rob_uop_2_2_pdst = {_RANDOM[11'h370][31], _RANDOM[11'h371][5:0]};	// rob.scala:310:28
        rob_uop_2_2_stale_pdst = _RANDOM[11'h372][10:4];	// rob.scala:310:28
        rob_uop_2_2_is_fencei = _RANDOM[11'h374][22];	// rob.scala:310:28
        rob_uop_2_2_uses_ldq = _RANDOM[11'h374][24];	// rob.scala:310:28
        rob_uop_2_2_uses_stq = _RANDOM[11'h374][25];	// rob.scala:310:28
        rob_uop_2_2_is_sys_pc2epc = _RANDOM[11'h374][26];	// rob.scala:310:28
        rob_uop_2_2_flush_on_commit = _RANDOM[11'h374][28];	// rob.scala:310:28
        rob_uop_2_2_ldst = {_RANDOM[11'h374][31:30], _RANDOM[11'h375][3:0]};	// rob.scala:310:28
        rob_uop_2_2_ldst_val = _RANDOM[11'h375][22];	// rob.scala:310:28
        rob_uop_2_2_dst_rtype = _RANDOM[11'h375][24:23];	// rob.scala:310:28
        rob_uop_2_2_fp_val = _RANDOM[11'h375][30];	// rob.scala:310:28
        rob_uop_2_3_uopc = _RANDOM[11'h376][15:9];	// rob.scala:310:28
        rob_uop_2_3_is_rvc = _RANDOM[11'h378][16];	// rob.scala:310:28
        rob_uop_2_3_br_mask = _RANDOM[11'h37B][20:5];	// rob.scala:310:28
        rob_uop_2_3_ftq_idx = _RANDOM[11'h37B][29:25];	// rob.scala:310:28
        rob_uop_2_3_edge_inst = _RANDOM[11'h37B][30];	// rob.scala:310:28
        rob_uop_2_3_pc_lob = {_RANDOM[11'h37B][31], _RANDOM[11'h37C][4:0]};	// rob.scala:310:28
        rob_uop_2_3_pdst = _RANDOM[11'h37D][31:25];	// rob.scala:310:28
        rob_uop_2_3_stale_pdst = {_RANDOM[11'h37E][31:30], _RANDOM[11'h37F][4:0]};	// rob.scala:310:28
        rob_uop_2_3_is_fencei = _RANDOM[11'h381][16];	// rob.scala:310:28
        rob_uop_2_3_uses_ldq = _RANDOM[11'h381][18];	// rob.scala:310:28
        rob_uop_2_3_uses_stq = _RANDOM[11'h381][19];	// rob.scala:310:28
        rob_uop_2_3_is_sys_pc2epc = _RANDOM[11'h381][20];	// rob.scala:310:28
        rob_uop_2_3_flush_on_commit = _RANDOM[11'h381][22];	// rob.scala:310:28
        rob_uop_2_3_ldst = _RANDOM[11'h381][29:24];	// rob.scala:310:28
        rob_uop_2_3_ldst_val = _RANDOM[11'h382][16];	// rob.scala:310:28
        rob_uop_2_3_dst_rtype = _RANDOM[11'h382][18:17];	// rob.scala:310:28
        rob_uop_2_3_fp_val = _RANDOM[11'h382][24];	// rob.scala:310:28
        rob_uop_2_4_uopc = _RANDOM[11'h383][9:3];	// rob.scala:310:28
        rob_uop_2_4_is_rvc = _RANDOM[11'h385][10];	// rob.scala:310:28
        rob_uop_2_4_br_mask = {_RANDOM[11'h387][31], _RANDOM[11'h388][14:0]};	// rob.scala:310:28
        rob_uop_2_4_ftq_idx = _RANDOM[11'h388][23:19];	// rob.scala:310:28
        rob_uop_2_4_edge_inst = _RANDOM[11'h388][24];	// rob.scala:310:28
        rob_uop_2_4_pc_lob = _RANDOM[11'h388][30:25];	// rob.scala:310:28
        rob_uop_2_4_pdst = _RANDOM[11'h38A][25:19];	// rob.scala:310:28
        rob_uop_2_4_stale_pdst = _RANDOM[11'h38B][30:24];	// rob.scala:310:28
        rob_uop_2_4_is_fencei = _RANDOM[11'h38E][10];	// rob.scala:310:28
        rob_uop_2_4_uses_ldq = _RANDOM[11'h38E][12];	// rob.scala:310:28
        rob_uop_2_4_uses_stq = _RANDOM[11'h38E][13];	// rob.scala:310:28
        rob_uop_2_4_is_sys_pc2epc = _RANDOM[11'h38E][14];	// rob.scala:310:28
        rob_uop_2_4_flush_on_commit = _RANDOM[11'h38E][16];	// rob.scala:310:28
        rob_uop_2_4_ldst = _RANDOM[11'h38E][23:18];	// rob.scala:310:28
        rob_uop_2_4_ldst_val = _RANDOM[11'h38F][10];	// rob.scala:310:28
        rob_uop_2_4_dst_rtype = _RANDOM[11'h38F][12:11];	// rob.scala:310:28
        rob_uop_2_4_fp_val = _RANDOM[11'h38F][18];	// rob.scala:310:28
        rob_uop_2_5_uopc = {_RANDOM[11'h38F][31:29], _RANDOM[11'h390][3:0]};	// rob.scala:310:28
        rob_uop_2_5_is_rvc = _RANDOM[11'h392][4];	// rob.scala:310:28
        rob_uop_2_5_br_mask = {_RANDOM[11'h394][31:25], _RANDOM[11'h395][8:0]};	// rob.scala:310:28
        rob_uop_2_5_ftq_idx = _RANDOM[11'h395][17:13];	// rob.scala:310:28
        rob_uop_2_5_edge_inst = _RANDOM[11'h395][18];	// rob.scala:310:28
        rob_uop_2_5_pc_lob = _RANDOM[11'h395][24:19];	// rob.scala:310:28
        rob_uop_2_5_pdst = _RANDOM[11'h397][19:13];	// rob.scala:310:28
        rob_uop_2_5_stale_pdst = _RANDOM[11'h398][24:18];	// rob.scala:310:28
        rob_uop_2_5_is_fencei = _RANDOM[11'h39B][4];	// rob.scala:310:28
        rob_uop_2_5_uses_ldq = _RANDOM[11'h39B][6];	// rob.scala:310:28
        rob_uop_2_5_uses_stq = _RANDOM[11'h39B][7];	// rob.scala:310:28
        rob_uop_2_5_is_sys_pc2epc = _RANDOM[11'h39B][8];	// rob.scala:310:28
        rob_uop_2_5_flush_on_commit = _RANDOM[11'h39B][10];	// rob.scala:310:28
        rob_uop_2_5_ldst = _RANDOM[11'h39B][17:12];	// rob.scala:310:28
        rob_uop_2_5_ldst_val = _RANDOM[11'h39C][4];	// rob.scala:310:28
        rob_uop_2_5_dst_rtype = _RANDOM[11'h39C][6:5];	// rob.scala:310:28
        rob_uop_2_5_fp_val = _RANDOM[11'h39C][12];	// rob.scala:310:28
        rob_uop_2_6_uopc = _RANDOM[11'h39C][29:23];	// rob.scala:310:28
        rob_uop_2_6_is_rvc = _RANDOM[11'h39E][30];	// rob.scala:310:28
        rob_uop_2_6_br_mask = {_RANDOM[11'h3A1][31:19], _RANDOM[11'h3A2][2:0]};	// rob.scala:310:28
        rob_uop_2_6_ftq_idx = _RANDOM[11'h3A2][11:7];	// rob.scala:310:28
        rob_uop_2_6_edge_inst = _RANDOM[11'h3A2][12];	// rob.scala:310:28
        rob_uop_2_6_pc_lob = _RANDOM[11'h3A2][18:13];	// rob.scala:310:28
        rob_uop_2_6_pdst = _RANDOM[11'h3A4][13:7];	// rob.scala:310:28
        rob_uop_2_6_stale_pdst = _RANDOM[11'h3A5][18:12];	// rob.scala:310:28
        rob_uop_2_6_is_fencei = _RANDOM[11'h3A7][30];	// rob.scala:310:28
        rob_uop_2_6_uses_ldq = _RANDOM[11'h3A8][0];	// rob.scala:310:28
        rob_uop_2_6_uses_stq = _RANDOM[11'h3A8][1];	// rob.scala:310:28
        rob_uop_2_6_is_sys_pc2epc = _RANDOM[11'h3A8][2];	// rob.scala:310:28
        rob_uop_2_6_flush_on_commit = _RANDOM[11'h3A8][4];	// rob.scala:310:28
        rob_uop_2_6_ldst = _RANDOM[11'h3A8][11:6];	// rob.scala:310:28
        rob_uop_2_6_ldst_val = _RANDOM[11'h3A8][30];	// rob.scala:310:28
        rob_uop_2_6_dst_rtype = {_RANDOM[11'h3A8][31], _RANDOM[11'h3A9][0]};	// rob.scala:310:28
        rob_uop_2_6_fp_val = _RANDOM[11'h3A9][6];	// rob.scala:310:28
        rob_uop_2_7_uopc = _RANDOM[11'h3A9][23:17];	// rob.scala:310:28
        rob_uop_2_7_is_rvc = _RANDOM[11'h3AB][24];	// rob.scala:310:28
        rob_uop_2_7_br_mask = _RANDOM[11'h3AE][28:13];	// rob.scala:310:28
        rob_uop_2_7_ftq_idx = _RANDOM[11'h3AF][5:1];	// rob.scala:310:28
        rob_uop_2_7_edge_inst = _RANDOM[11'h3AF][6];	// rob.scala:310:28
        rob_uop_2_7_pc_lob = _RANDOM[11'h3AF][12:7];	// rob.scala:310:28
        rob_uop_2_7_pdst = _RANDOM[11'h3B1][7:1];	// rob.scala:310:28
        rob_uop_2_7_stale_pdst = _RANDOM[11'h3B2][12:6];	// rob.scala:310:28
        rob_uop_2_7_is_fencei = _RANDOM[11'h3B4][24];	// rob.scala:310:28
        rob_uop_2_7_uses_ldq = _RANDOM[11'h3B4][26];	// rob.scala:310:28
        rob_uop_2_7_uses_stq = _RANDOM[11'h3B4][27];	// rob.scala:310:28
        rob_uop_2_7_is_sys_pc2epc = _RANDOM[11'h3B4][28];	// rob.scala:310:28
        rob_uop_2_7_flush_on_commit = _RANDOM[11'h3B4][30];	// rob.scala:310:28
        rob_uop_2_7_ldst = _RANDOM[11'h3B5][5:0];	// rob.scala:310:28
        rob_uop_2_7_ldst_val = _RANDOM[11'h3B5][24];	// rob.scala:310:28
        rob_uop_2_7_dst_rtype = _RANDOM[11'h3B5][26:25];	// rob.scala:310:28
        rob_uop_2_7_fp_val = _RANDOM[11'h3B6][0];	// rob.scala:310:28
        rob_uop_2_8_uopc = _RANDOM[11'h3B6][17:11];	// rob.scala:310:28
        rob_uop_2_8_is_rvc = _RANDOM[11'h3B8][18];	// rob.scala:310:28
        rob_uop_2_8_br_mask = _RANDOM[11'h3BB][22:7];	// rob.scala:310:28
        rob_uop_2_8_ftq_idx = _RANDOM[11'h3BB][31:27];	// rob.scala:310:28
        rob_uop_2_8_edge_inst = _RANDOM[11'h3BC][0];	// rob.scala:310:28
        rob_uop_2_8_pc_lob = _RANDOM[11'h3BC][6:1];	// rob.scala:310:28
        rob_uop_2_8_pdst = {_RANDOM[11'h3BD][31:27], _RANDOM[11'h3BE][1:0]};	// rob.scala:310:28
        rob_uop_2_8_stale_pdst = _RANDOM[11'h3BF][6:0];	// rob.scala:310:28
        rob_uop_2_8_is_fencei = _RANDOM[11'h3C1][18];	// rob.scala:310:28
        rob_uop_2_8_uses_ldq = _RANDOM[11'h3C1][20];	// rob.scala:310:28
        rob_uop_2_8_uses_stq = _RANDOM[11'h3C1][21];	// rob.scala:310:28
        rob_uop_2_8_is_sys_pc2epc = _RANDOM[11'h3C1][22];	// rob.scala:310:28
        rob_uop_2_8_flush_on_commit = _RANDOM[11'h3C1][24];	// rob.scala:310:28
        rob_uop_2_8_ldst = _RANDOM[11'h3C1][31:26];	// rob.scala:310:28
        rob_uop_2_8_ldst_val = _RANDOM[11'h3C2][18];	// rob.scala:310:28
        rob_uop_2_8_dst_rtype = _RANDOM[11'h3C2][20:19];	// rob.scala:310:28
        rob_uop_2_8_fp_val = _RANDOM[11'h3C2][26];	// rob.scala:310:28
        rob_uop_2_9_uopc = _RANDOM[11'h3C3][11:5];	// rob.scala:310:28
        rob_uop_2_9_is_rvc = _RANDOM[11'h3C5][12];	// rob.scala:310:28
        rob_uop_2_9_br_mask = _RANDOM[11'h3C8][16:1];	// rob.scala:310:28
        rob_uop_2_9_ftq_idx = _RANDOM[11'h3C8][25:21];	// rob.scala:310:28
        rob_uop_2_9_edge_inst = _RANDOM[11'h3C8][26];	// rob.scala:310:28
        rob_uop_2_9_pc_lob = {_RANDOM[11'h3C8][31:27], _RANDOM[11'h3C9][0]};	// rob.scala:310:28
        rob_uop_2_9_pdst = _RANDOM[11'h3CA][27:21];	// rob.scala:310:28
        rob_uop_2_9_stale_pdst = {_RANDOM[11'h3CB][31:26], _RANDOM[11'h3CC][0]};	// rob.scala:310:28
        rob_uop_2_9_is_fencei = _RANDOM[11'h3CE][12];	// rob.scala:310:28
        rob_uop_2_9_uses_ldq = _RANDOM[11'h3CE][14];	// rob.scala:310:28
        rob_uop_2_9_uses_stq = _RANDOM[11'h3CE][15];	// rob.scala:310:28
        rob_uop_2_9_is_sys_pc2epc = _RANDOM[11'h3CE][16];	// rob.scala:310:28
        rob_uop_2_9_flush_on_commit = _RANDOM[11'h3CE][18];	// rob.scala:310:28
        rob_uop_2_9_ldst = _RANDOM[11'h3CE][25:20];	// rob.scala:310:28
        rob_uop_2_9_ldst_val = _RANDOM[11'h3CF][12];	// rob.scala:310:28
        rob_uop_2_9_dst_rtype = _RANDOM[11'h3CF][14:13];	// rob.scala:310:28
        rob_uop_2_9_fp_val = _RANDOM[11'h3CF][20];	// rob.scala:310:28
        rob_uop_2_10_uopc = {_RANDOM[11'h3CF][31], _RANDOM[11'h3D0][5:0]};	// rob.scala:310:28
        rob_uop_2_10_is_rvc = _RANDOM[11'h3D2][6];	// rob.scala:310:28
        rob_uop_2_10_br_mask = {_RANDOM[11'h3D4][31:27], _RANDOM[11'h3D5][10:0]};	// rob.scala:310:28
        rob_uop_2_10_ftq_idx = _RANDOM[11'h3D5][19:15];	// rob.scala:310:28
        rob_uop_2_10_edge_inst = _RANDOM[11'h3D5][20];	// rob.scala:310:28
        rob_uop_2_10_pc_lob = _RANDOM[11'h3D5][26:21];	// rob.scala:310:28
        rob_uop_2_10_pdst = _RANDOM[11'h3D7][21:15];	// rob.scala:310:28
        rob_uop_2_10_stale_pdst = _RANDOM[11'h3D8][26:20];	// rob.scala:310:28
        rob_uop_2_10_is_fencei = _RANDOM[11'h3DB][6];	// rob.scala:310:28
        rob_uop_2_10_uses_ldq = _RANDOM[11'h3DB][8];	// rob.scala:310:28
        rob_uop_2_10_uses_stq = _RANDOM[11'h3DB][9];	// rob.scala:310:28
        rob_uop_2_10_is_sys_pc2epc = _RANDOM[11'h3DB][10];	// rob.scala:310:28
        rob_uop_2_10_flush_on_commit = _RANDOM[11'h3DB][12];	// rob.scala:310:28
        rob_uop_2_10_ldst = _RANDOM[11'h3DB][19:14];	// rob.scala:310:28
        rob_uop_2_10_ldst_val = _RANDOM[11'h3DC][6];	// rob.scala:310:28
        rob_uop_2_10_dst_rtype = _RANDOM[11'h3DC][8:7];	// rob.scala:310:28
        rob_uop_2_10_fp_val = _RANDOM[11'h3DC][14];	// rob.scala:310:28
        rob_uop_2_11_uopc = _RANDOM[11'h3DC][31:25];	// rob.scala:310:28
        rob_uop_2_11_is_rvc = _RANDOM[11'h3DF][0];	// rob.scala:310:28
        rob_uop_2_11_br_mask = {_RANDOM[11'h3E1][31:21], _RANDOM[11'h3E2][4:0]};	// rob.scala:310:28
        rob_uop_2_11_ftq_idx = _RANDOM[11'h3E2][13:9];	// rob.scala:310:28
        rob_uop_2_11_edge_inst = _RANDOM[11'h3E2][14];	// rob.scala:310:28
        rob_uop_2_11_pc_lob = _RANDOM[11'h3E2][20:15];	// rob.scala:310:28
        rob_uop_2_11_pdst = _RANDOM[11'h3E4][15:9];	// rob.scala:310:28
        rob_uop_2_11_stale_pdst = _RANDOM[11'h3E5][20:14];	// rob.scala:310:28
        rob_uop_2_11_is_fencei = _RANDOM[11'h3E8][0];	// rob.scala:310:28
        rob_uop_2_11_uses_ldq = _RANDOM[11'h3E8][2];	// rob.scala:310:28
        rob_uop_2_11_uses_stq = _RANDOM[11'h3E8][3];	// rob.scala:310:28
        rob_uop_2_11_is_sys_pc2epc = _RANDOM[11'h3E8][4];	// rob.scala:310:28
        rob_uop_2_11_flush_on_commit = _RANDOM[11'h3E8][6];	// rob.scala:310:28
        rob_uop_2_11_ldst = _RANDOM[11'h3E8][13:8];	// rob.scala:310:28
        rob_uop_2_11_ldst_val = _RANDOM[11'h3E9][0];	// rob.scala:310:28
        rob_uop_2_11_dst_rtype = _RANDOM[11'h3E9][2:1];	// rob.scala:310:28
        rob_uop_2_11_fp_val = _RANDOM[11'h3E9][8];	// rob.scala:310:28
        rob_uop_2_12_uopc = _RANDOM[11'h3E9][25:19];	// rob.scala:310:28
        rob_uop_2_12_is_rvc = _RANDOM[11'h3EB][26];	// rob.scala:310:28
        rob_uop_2_12_br_mask = _RANDOM[11'h3EE][30:15];	// rob.scala:310:28
        rob_uop_2_12_ftq_idx = _RANDOM[11'h3EF][7:3];	// rob.scala:310:28
        rob_uop_2_12_edge_inst = _RANDOM[11'h3EF][8];	// rob.scala:310:28
        rob_uop_2_12_pc_lob = _RANDOM[11'h3EF][14:9];	// rob.scala:310:28
        rob_uop_2_12_pdst = _RANDOM[11'h3F1][9:3];	// rob.scala:310:28
        rob_uop_2_12_stale_pdst = _RANDOM[11'h3F2][14:8];	// rob.scala:310:28
        rob_uop_2_12_is_fencei = _RANDOM[11'h3F4][26];	// rob.scala:310:28
        rob_uop_2_12_uses_ldq = _RANDOM[11'h3F4][28];	// rob.scala:310:28
        rob_uop_2_12_uses_stq = _RANDOM[11'h3F4][29];	// rob.scala:310:28
        rob_uop_2_12_is_sys_pc2epc = _RANDOM[11'h3F4][30];	// rob.scala:310:28
        rob_uop_2_12_flush_on_commit = _RANDOM[11'h3F5][0];	// rob.scala:310:28
        rob_uop_2_12_ldst = _RANDOM[11'h3F5][7:2];	// rob.scala:310:28
        rob_uop_2_12_ldst_val = _RANDOM[11'h3F5][26];	// rob.scala:310:28
        rob_uop_2_12_dst_rtype = _RANDOM[11'h3F5][28:27];	// rob.scala:310:28
        rob_uop_2_12_fp_val = _RANDOM[11'h3F6][2];	// rob.scala:310:28
        rob_uop_2_13_uopc = _RANDOM[11'h3F6][19:13];	// rob.scala:310:28
        rob_uop_2_13_is_rvc = _RANDOM[11'h3F8][20];	// rob.scala:310:28
        rob_uop_2_13_br_mask = _RANDOM[11'h3FB][24:9];	// rob.scala:310:28
        rob_uop_2_13_ftq_idx = {_RANDOM[11'h3FB][31:29], _RANDOM[11'h3FC][1:0]};	// rob.scala:310:28
        rob_uop_2_13_edge_inst = _RANDOM[11'h3FC][2];	// rob.scala:310:28
        rob_uop_2_13_pc_lob = _RANDOM[11'h3FC][8:3];	// rob.scala:310:28
        rob_uop_2_13_pdst = {_RANDOM[11'h3FD][31:29], _RANDOM[11'h3FE][3:0]};	// rob.scala:310:28
        rob_uop_2_13_stale_pdst = _RANDOM[11'h3FF][8:2];	// rob.scala:310:28
        rob_uop_2_13_is_fencei = _RANDOM[11'h401][20];	// rob.scala:310:28
        rob_uop_2_13_uses_ldq = _RANDOM[11'h401][22];	// rob.scala:310:28
        rob_uop_2_13_uses_stq = _RANDOM[11'h401][23];	// rob.scala:310:28
        rob_uop_2_13_is_sys_pc2epc = _RANDOM[11'h401][24];	// rob.scala:310:28
        rob_uop_2_13_flush_on_commit = _RANDOM[11'h401][26];	// rob.scala:310:28
        rob_uop_2_13_ldst = {_RANDOM[11'h401][31:28], _RANDOM[11'h402][1:0]};	// rob.scala:310:28
        rob_uop_2_13_ldst_val = _RANDOM[11'h402][20];	// rob.scala:310:28
        rob_uop_2_13_dst_rtype = _RANDOM[11'h402][22:21];	// rob.scala:310:28
        rob_uop_2_13_fp_val = _RANDOM[11'h402][28];	// rob.scala:310:28
        rob_uop_2_14_uopc = _RANDOM[11'h403][13:7];	// rob.scala:310:28
        rob_uop_2_14_is_rvc = _RANDOM[11'h405][14];	// rob.scala:310:28
        rob_uop_2_14_br_mask = _RANDOM[11'h408][18:3];	// rob.scala:310:28
        rob_uop_2_14_ftq_idx = _RANDOM[11'h408][27:23];	// rob.scala:310:28
        rob_uop_2_14_edge_inst = _RANDOM[11'h408][28];	// rob.scala:310:28
        rob_uop_2_14_pc_lob = {_RANDOM[11'h408][31:29], _RANDOM[11'h409][2:0]};	// rob.scala:310:28
        rob_uop_2_14_pdst = _RANDOM[11'h40A][29:23];	// rob.scala:310:28
        rob_uop_2_14_stale_pdst = {_RANDOM[11'h40B][31:28], _RANDOM[11'h40C][2:0]};	// rob.scala:310:28
        rob_uop_2_14_is_fencei = _RANDOM[11'h40E][14];	// rob.scala:310:28
        rob_uop_2_14_uses_ldq = _RANDOM[11'h40E][16];	// rob.scala:310:28
        rob_uop_2_14_uses_stq = _RANDOM[11'h40E][17];	// rob.scala:310:28
        rob_uop_2_14_is_sys_pc2epc = _RANDOM[11'h40E][18];	// rob.scala:310:28
        rob_uop_2_14_flush_on_commit = _RANDOM[11'h40E][20];	// rob.scala:310:28
        rob_uop_2_14_ldst = _RANDOM[11'h40E][27:22];	// rob.scala:310:28
        rob_uop_2_14_ldst_val = _RANDOM[11'h40F][14];	// rob.scala:310:28
        rob_uop_2_14_dst_rtype = _RANDOM[11'h40F][16:15];	// rob.scala:310:28
        rob_uop_2_14_fp_val = _RANDOM[11'h40F][22];	// rob.scala:310:28
        rob_uop_2_15_uopc = _RANDOM[11'h410][7:1];	// rob.scala:310:28
        rob_uop_2_15_is_rvc = _RANDOM[11'h412][8];	// rob.scala:310:28
        rob_uop_2_15_br_mask = {_RANDOM[11'h414][31:29], _RANDOM[11'h415][12:0]};	// rob.scala:310:28
        rob_uop_2_15_ftq_idx = _RANDOM[11'h415][21:17];	// rob.scala:310:28
        rob_uop_2_15_edge_inst = _RANDOM[11'h415][22];	// rob.scala:310:28
        rob_uop_2_15_pc_lob = _RANDOM[11'h415][28:23];	// rob.scala:310:28
        rob_uop_2_15_pdst = _RANDOM[11'h417][23:17];	// rob.scala:310:28
        rob_uop_2_15_stale_pdst = _RANDOM[11'h418][28:22];	// rob.scala:310:28
        rob_uop_2_15_is_fencei = _RANDOM[11'h41B][8];	// rob.scala:310:28
        rob_uop_2_15_uses_ldq = _RANDOM[11'h41B][10];	// rob.scala:310:28
        rob_uop_2_15_uses_stq = _RANDOM[11'h41B][11];	// rob.scala:310:28
        rob_uop_2_15_is_sys_pc2epc = _RANDOM[11'h41B][12];	// rob.scala:310:28
        rob_uop_2_15_flush_on_commit = _RANDOM[11'h41B][14];	// rob.scala:310:28
        rob_uop_2_15_ldst = _RANDOM[11'h41B][21:16];	// rob.scala:310:28
        rob_uop_2_15_ldst_val = _RANDOM[11'h41C][8];	// rob.scala:310:28
        rob_uop_2_15_dst_rtype = _RANDOM[11'h41C][10:9];	// rob.scala:310:28
        rob_uop_2_15_fp_val = _RANDOM[11'h41C][16];	// rob.scala:310:28
        rob_uop_2_16_uopc = {_RANDOM[11'h41C][31:27], _RANDOM[11'h41D][1:0]};	// rob.scala:310:28
        rob_uop_2_16_is_rvc = _RANDOM[11'h41F][2];	// rob.scala:310:28
        rob_uop_2_16_br_mask = {_RANDOM[11'h421][31:23], _RANDOM[11'h422][6:0]};	// rob.scala:310:28
        rob_uop_2_16_ftq_idx = _RANDOM[11'h422][15:11];	// rob.scala:310:28
        rob_uop_2_16_edge_inst = _RANDOM[11'h422][16];	// rob.scala:310:28
        rob_uop_2_16_pc_lob = _RANDOM[11'h422][22:17];	// rob.scala:310:28
        rob_uop_2_16_pdst = _RANDOM[11'h424][17:11];	// rob.scala:310:28
        rob_uop_2_16_stale_pdst = _RANDOM[11'h425][22:16];	// rob.scala:310:28
        rob_uop_2_16_is_fencei = _RANDOM[11'h428][2];	// rob.scala:310:28
        rob_uop_2_16_uses_ldq = _RANDOM[11'h428][4];	// rob.scala:310:28
        rob_uop_2_16_uses_stq = _RANDOM[11'h428][5];	// rob.scala:310:28
        rob_uop_2_16_is_sys_pc2epc = _RANDOM[11'h428][6];	// rob.scala:310:28
        rob_uop_2_16_flush_on_commit = _RANDOM[11'h428][8];	// rob.scala:310:28
        rob_uop_2_16_ldst = _RANDOM[11'h428][15:10];	// rob.scala:310:28
        rob_uop_2_16_ldst_val = _RANDOM[11'h429][2];	// rob.scala:310:28
        rob_uop_2_16_dst_rtype = _RANDOM[11'h429][4:3];	// rob.scala:310:28
        rob_uop_2_16_fp_val = _RANDOM[11'h429][10];	// rob.scala:310:28
        rob_uop_2_17_uopc = _RANDOM[11'h429][27:21];	// rob.scala:310:28
        rob_uop_2_17_is_rvc = _RANDOM[11'h42B][28];	// rob.scala:310:28
        rob_uop_2_17_br_mask = {_RANDOM[11'h42E][31:17], _RANDOM[11'h42F][0]};	// rob.scala:310:28
        rob_uop_2_17_ftq_idx = _RANDOM[11'h42F][9:5];	// rob.scala:310:28
        rob_uop_2_17_edge_inst = _RANDOM[11'h42F][10];	// rob.scala:310:28
        rob_uop_2_17_pc_lob = _RANDOM[11'h42F][16:11];	// rob.scala:310:28
        rob_uop_2_17_pdst = _RANDOM[11'h431][11:5];	// rob.scala:310:28
        rob_uop_2_17_stale_pdst = _RANDOM[11'h432][16:10];	// rob.scala:310:28
        rob_uop_2_17_is_fencei = _RANDOM[11'h434][28];	// rob.scala:310:28
        rob_uop_2_17_uses_ldq = _RANDOM[11'h434][30];	// rob.scala:310:28
        rob_uop_2_17_uses_stq = _RANDOM[11'h434][31];	// rob.scala:310:28
        rob_uop_2_17_is_sys_pc2epc = _RANDOM[11'h435][0];	// rob.scala:310:28
        rob_uop_2_17_flush_on_commit = _RANDOM[11'h435][2];	// rob.scala:310:28
        rob_uop_2_17_ldst = _RANDOM[11'h435][9:4];	// rob.scala:310:28
        rob_uop_2_17_ldst_val = _RANDOM[11'h435][28];	// rob.scala:310:28
        rob_uop_2_17_dst_rtype = _RANDOM[11'h435][30:29];	// rob.scala:310:28
        rob_uop_2_17_fp_val = _RANDOM[11'h436][4];	// rob.scala:310:28
        rob_uop_2_18_uopc = _RANDOM[11'h436][21:15];	// rob.scala:310:28
        rob_uop_2_18_is_rvc = _RANDOM[11'h438][22];	// rob.scala:310:28
        rob_uop_2_18_br_mask = _RANDOM[11'h43B][26:11];	// rob.scala:310:28
        rob_uop_2_18_ftq_idx = {_RANDOM[11'h43B][31], _RANDOM[11'h43C][3:0]};	// rob.scala:310:28
        rob_uop_2_18_edge_inst = _RANDOM[11'h43C][4];	// rob.scala:310:28
        rob_uop_2_18_pc_lob = _RANDOM[11'h43C][10:5];	// rob.scala:310:28
        rob_uop_2_18_pdst = {_RANDOM[11'h43D][31], _RANDOM[11'h43E][5:0]};	// rob.scala:310:28
        rob_uop_2_18_stale_pdst = _RANDOM[11'h43F][10:4];	// rob.scala:310:28
        rob_uop_2_18_is_fencei = _RANDOM[11'h441][22];	// rob.scala:310:28
        rob_uop_2_18_uses_ldq = _RANDOM[11'h441][24];	// rob.scala:310:28
        rob_uop_2_18_uses_stq = _RANDOM[11'h441][25];	// rob.scala:310:28
        rob_uop_2_18_is_sys_pc2epc = _RANDOM[11'h441][26];	// rob.scala:310:28
        rob_uop_2_18_flush_on_commit = _RANDOM[11'h441][28];	// rob.scala:310:28
        rob_uop_2_18_ldst = {_RANDOM[11'h441][31:30], _RANDOM[11'h442][3:0]};	// rob.scala:310:28
        rob_uop_2_18_ldst_val = _RANDOM[11'h442][22];	// rob.scala:310:28
        rob_uop_2_18_dst_rtype = _RANDOM[11'h442][24:23];	// rob.scala:310:28
        rob_uop_2_18_fp_val = _RANDOM[11'h442][30];	// rob.scala:310:28
        rob_uop_2_19_uopc = _RANDOM[11'h443][15:9];	// rob.scala:310:28
        rob_uop_2_19_is_rvc = _RANDOM[11'h445][16];	// rob.scala:310:28
        rob_uop_2_19_br_mask = _RANDOM[11'h448][20:5];	// rob.scala:310:28
        rob_uop_2_19_ftq_idx = _RANDOM[11'h448][29:25];	// rob.scala:310:28
        rob_uop_2_19_edge_inst = _RANDOM[11'h448][30];	// rob.scala:310:28
        rob_uop_2_19_pc_lob = {_RANDOM[11'h448][31], _RANDOM[11'h449][4:0]};	// rob.scala:310:28
        rob_uop_2_19_pdst = _RANDOM[11'h44A][31:25];	// rob.scala:310:28
        rob_uop_2_19_stale_pdst = {_RANDOM[11'h44B][31:30], _RANDOM[11'h44C][4:0]};	// rob.scala:310:28
        rob_uop_2_19_is_fencei = _RANDOM[11'h44E][16];	// rob.scala:310:28
        rob_uop_2_19_uses_ldq = _RANDOM[11'h44E][18];	// rob.scala:310:28
        rob_uop_2_19_uses_stq = _RANDOM[11'h44E][19];	// rob.scala:310:28
        rob_uop_2_19_is_sys_pc2epc = _RANDOM[11'h44E][20];	// rob.scala:310:28
        rob_uop_2_19_flush_on_commit = _RANDOM[11'h44E][22];	// rob.scala:310:28
        rob_uop_2_19_ldst = _RANDOM[11'h44E][29:24];	// rob.scala:310:28
        rob_uop_2_19_ldst_val = _RANDOM[11'h44F][16];	// rob.scala:310:28
        rob_uop_2_19_dst_rtype = _RANDOM[11'h44F][18:17];	// rob.scala:310:28
        rob_uop_2_19_fp_val = _RANDOM[11'h44F][24];	// rob.scala:310:28
        rob_uop_2_20_uopc = _RANDOM[11'h450][9:3];	// rob.scala:310:28
        rob_uop_2_20_is_rvc = _RANDOM[11'h452][10];	// rob.scala:310:28
        rob_uop_2_20_br_mask = {_RANDOM[11'h454][31], _RANDOM[11'h455][14:0]};	// rob.scala:310:28
        rob_uop_2_20_ftq_idx = _RANDOM[11'h455][23:19];	// rob.scala:310:28
        rob_uop_2_20_edge_inst = _RANDOM[11'h455][24];	// rob.scala:310:28
        rob_uop_2_20_pc_lob = _RANDOM[11'h455][30:25];	// rob.scala:310:28
        rob_uop_2_20_pdst = _RANDOM[11'h457][25:19];	// rob.scala:310:28
        rob_uop_2_20_stale_pdst = _RANDOM[11'h458][30:24];	// rob.scala:310:28
        rob_uop_2_20_is_fencei = _RANDOM[11'h45B][10];	// rob.scala:310:28
        rob_uop_2_20_uses_ldq = _RANDOM[11'h45B][12];	// rob.scala:310:28
        rob_uop_2_20_uses_stq = _RANDOM[11'h45B][13];	// rob.scala:310:28
        rob_uop_2_20_is_sys_pc2epc = _RANDOM[11'h45B][14];	// rob.scala:310:28
        rob_uop_2_20_flush_on_commit = _RANDOM[11'h45B][16];	// rob.scala:310:28
        rob_uop_2_20_ldst = _RANDOM[11'h45B][23:18];	// rob.scala:310:28
        rob_uop_2_20_ldst_val = _RANDOM[11'h45C][10];	// rob.scala:310:28
        rob_uop_2_20_dst_rtype = _RANDOM[11'h45C][12:11];	// rob.scala:310:28
        rob_uop_2_20_fp_val = _RANDOM[11'h45C][18];	// rob.scala:310:28
        rob_uop_2_21_uopc = {_RANDOM[11'h45C][31:29], _RANDOM[11'h45D][3:0]};	// rob.scala:310:28
        rob_uop_2_21_is_rvc = _RANDOM[11'h45F][4];	// rob.scala:310:28
        rob_uop_2_21_br_mask = {_RANDOM[11'h461][31:25], _RANDOM[11'h462][8:0]};	// rob.scala:310:28
        rob_uop_2_21_ftq_idx = _RANDOM[11'h462][17:13];	// rob.scala:310:28
        rob_uop_2_21_edge_inst = _RANDOM[11'h462][18];	// rob.scala:310:28
        rob_uop_2_21_pc_lob = _RANDOM[11'h462][24:19];	// rob.scala:310:28
        rob_uop_2_21_pdst = _RANDOM[11'h464][19:13];	// rob.scala:310:28
        rob_uop_2_21_stale_pdst = _RANDOM[11'h465][24:18];	// rob.scala:310:28
        rob_uop_2_21_is_fencei = _RANDOM[11'h468][4];	// rob.scala:310:28
        rob_uop_2_21_uses_ldq = _RANDOM[11'h468][6];	// rob.scala:310:28
        rob_uop_2_21_uses_stq = _RANDOM[11'h468][7];	// rob.scala:310:28
        rob_uop_2_21_is_sys_pc2epc = _RANDOM[11'h468][8];	// rob.scala:310:28
        rob_uop_2_21_flush_on_commit = _RANDOM[11'h468][10];	// rob.scala:310:28
        rob_uop_2_21_ldst = _RANDOM[11'h468][17:12];	// rob.scala:310:28
        rob_uop_2_21_ldst_val = _RANDOM[11'h469][4];	// rob.scala:310:28
        rob_uop_2_21_dst_rtype = _RANDOM[11'h469][6:5];	// rob.scala:310:28
        rob_uop_2_21_fp_val = _RANDOM[11'h469][12];	// rob.scala:310:28
        rob_uop_2_22_uopc = _RANDOM[11'h469][29:23];	// rob.scala:310:28
        rob_uop_2_22_is_rvc = _RANDOM[11'h46B][30];	// rob.scala:310:28
        rob_uop_2_22_br_mask = {_RANDOM[11'h46E][31:19], _RANDOM[11'h46F][2:0]};	// rob.scala:310:28
        rob_uop_2_22_ftq_idx = _RANDOM[11'h46F][11:7];	// rob.scala:310:28
        rob_uop_2_22_edge_inst = _RANDOM[11'h46F][12];	// rob.scala:310:28
        rob_uop_2_22_pc_lob = _RANDOM[11'h46F][18:13];	// rob.scala:310:28
        rob_uop_2_22_pdst = _RANDOM[11'h471][13:7];	// rob.scala:310:28
        rob_uop_2_22_stale_pdst = _RANDOM[11'h472][18:12];	// rob.scala:310:28
        rob_uop_2_22_is_fencei = _RANDOM[11'h474][30];	// rob.scala:310:28
        rob_uop_2_22_uses_ldq = _RANDOM[11'h475][0];	// rob.scala:310:28
        rob_uop_2_22_uses_stq = _RANDOM[11'h475][1];	// rob.scala:310:28
        rob_uop_2_22_is_sys_pc2epc = _RANDOM[11'h475][2];	// rob.scala:310:28
        rob_uop_2_22_flush_on_commit = _RANDOM[11'h475][4];	// rob.scala:310:28
        rob_uop_2_22_ldst = _RANDOM[11'h475][11:6];	// rob.scala:310:28
        rob_uop_2_22_ldst_val = _RANDOM[11'h475][30];	// rob.scala:310:28
        rob_uop_2_22_dst_rtype = {_RANDOM[11'h475][31], _RANDOM[11'h476][0]};	// rob.scala:310:28
        rob_uop_2_22_fp_val = _RANDOM[11'h476][6];	// rob.scala:310:28
        rob_uop_2_23_uopc = _RANDOM[11'h476][23:17];	// rob.scala:310:28
        rob_uop_2_23_is_rvc = _RANDOM[11'h478][24];	// rob.scala:310:28
        rob_uop_2_23_br_mask = _RANDOM[11'h47B][28:13];	// rob.scala:310:28
        rob_uop_2_23_ftq_idx = _RANDOM[11'h47C][5:1];	// rob.scala:310:28
        rob_uop_2_23_edge_inst = _RANDOM[11'h47C][6];	// rob.scala:310:28
        rob_uop_2_23_pc_lob = _RANDOM[11'h47C][12:7];	// rob.scala:310:28
        rob_uop_2_23_pdst = _RANDOM[11'h47E][7:1];	// rob.scala:310:28
        rob_uop_2_23_stale_pdst = _RANDOM[11'h47F][12:6];	// rob.scala:310:28
        rob_uop_2_23_is_fencei = _RANDOM[11'h481][24];	// rob.scala:310:28
        rob_uop_2_23_uses_ldq = _RANDOM[11'h481][26];	// rob.scala:310:28
        rob_uop_2_23_uses_stq = _RANDOM[11'h481][27];	// rob.scala:310:28
        rob_uop_2_23_is_sys_pc2epc = _RANDOM[11'h481][28];	// rob.scala:310:28
        rob_uop_2_23_flush_on_commit = _RANDOM[11'h481][30];	// rob.scala:310:28
        rob_uop_2_23_ldst = _RANDOM[11'h482][5:0];	// rob.scala:310:28
        rob_uop_2_23_ldst_val = _RANDOM[11'h482][24];	// rob.scala:310:28
        rob_uop_2_23_dst_rtype = _RANDOM[11'h482][26:25];	// rob.scala:310:28
        rob_uop_2_23_fp_val = _RANDOM[11'h483][0];	// rob.scala:310:28
        rob_uop_2_24_uopc = _RANDOM[11'h483][17:11];	// rob.scala:310:28
        rob_uop_2_24_is_rvc = _RANDOM[11'h485][18];	// rob.scala:310:28
        rob_uop_2_24_br_mask = _RANDOM[11'h488][22:7];	// rob.scala:310:28
        rob_uop_2_24_ftq_idx = _RANDOM[11'h488][31:27];	// rob.scala:310:28
        rob_uop_2_24_edge_inst = _RANDOM[11'h489][0];	// rob.scala:310:28
        rob_uop_2_24_pc_lob = _RANDOM[11'h489][6:1];	// rob.scala:310:28
        rob_uop_2_24_pdst = {_RANDOM[11'h48A][31:27], _RANDOM[11'h48B][1:0]};	// rob.scala:310:28
        rob_uop_2_24_stale_pdst = _RANDOM[11'h48C][6:0];	// rob.scala:310:28
        rob_uop_2_24_is_fencei = _RANDOM[11'h48E][18];	// rob.scala:310:28
        rob_uop_2_24_uses_ldq = _RANDOM[11'h48E][20];	// rob.scala:310:28
        rob_uop_2_24_uses_stq = _RANDOM[11'h48E][21];	// rob.scala:310:28
        rob_uop_2_24_is_sys_pc2epc = _RANDOM[11'h48E][22];	// rob.scala:310:28
        rob_uop_2_24_flush_on_commit = _RANDOM[11'h48E][24];	// rob.scala:310:28
        rob_uop_2_24_ldst = _RANDOM[11'h48E][31:26];	// rob.scala:310:28
        rob_uop_2_24_ldst_val = _RANDOM[11'h48F][18];	// rob.scala:310:28
        rob_uop_2_24_dst_rtype = _RANDOM[11'h48F][20:19];	// rob.scala:310:28
        rob_uop_2_24_fp_val = _RANDOM[11'h48F][26];	// rob.scala:310:28
        rob_uop_2_25_uopc = _RANDOM[11'h490][11:5];	// rob.scala:310:28
        rob_uop_2_25_is_rvc = _RANDOM[11'h492][12];	// rob.scala:310:28
        rob_uop_2_25_br_mask = _RANDOM[11'h495][16:1];	// rob.scala:310:28
        rob_uop_2_25_ftq_idx = _RANDOM[11'h495][25:21];	// rob.scala:310:28
        rob_uop_2_25_edge_inst = _RANDOM[11'h495][26];	// rob.scala:310:28
        rob_uop_2_25_pc_lob = {_RANDOM[11'h495][31:27], _RANDOM[11'h496][0]};	// rob.scala:310:28
        rob_uop_2_25_pdst = _RANDOM[11'h497][27:21];	// rob.scala:310:28
        rob_uop_2_25_stale_pdst = {_RANDOM[11'h498][31:26], _RANDOM[11'h499][0]};	// rob.scala:310:28
        rob_uop_2_25_is_fencei = _RANDOM[11'h49B][12];	// rob.scala:310:28
        rob_uop_2_25_uses_ldq = _RANDOM[11'h49B][14];	// rob.scala:310:28
        rob_uop_2_25_uses_stq = _RANDOM[11'h49B][15];	// rob.scala:310:28
        rob_uop_2_25_is_sys_pc2epc = _RANDOM[11'h49B][16];	// rob.scala:310:28
        rob_uop_2_25_flush_on_commit = _RANDOM[11'h49B][18];	// rob.scala:310:28
        rob_uop_2_25_ldst = _RANDOM[11'h49B][25:20];	// rob.scala:310:28
        rob_uop_2_25_ldst_val = _RANDOM[11'h49C][12];	// rob.scala:310:28
        rob_uop_2_25_dst_rtype = _RANDOM[11'h49C][14:13];	// rob.scala:310:28
        rob_uop_2_25_fp_val = _RANDOM[11'h49C][20];	// rob.scala:310:28
        rob_uop_2_26_uopc = {_RANDOM[11'h49C][31], _RANDOM[11'h49D][5:0]};	// rob.scala:310:28
        rob_uop_2_26_is_rvc = _RANDOM[11'h49F][6];	// rob.scala:310:28
        rob_uop_2_26_br_mask = {_RANDOM[11'h4A1][31:27], _RANDOM[11'h4A2][10:0]};	// rob.scala:310:28
        rob_uop_2_26_ftq_idx = _RANDOM[11'h4A2][19:15];	// rob.scala:310:28
        rob_uop_2_26_edge_inst = _RANDOM[11'h4A2][20];	// rob.scala:310:28
        rob_uop_2_26_pc_lob = _RANDOM[11'h4A2][26:21];	// rob.scala:310:28
        rob_uop_2_26_pdst = _RANDOM[11'h4A4][21:15];	// rob.scala:310:28
        rob_uop_2_26_stale_pdst = _RANDOM[11'h4A5][26:20];	// rob.scala:310:28
        rob_uop_2_26_is_fencei = _RANDOM[11'h4A8][6];	// rob.scala:310:28
        rob_uop_2_26_uses_ldq = _RANDOM[11'h4A8][8];	// rob.scala:310:28
        rob_uop_2_26_uses_stq = _RANDOM[11'h4A8][9];	// rob.scala:310:28
        rob_uop_2_26_is_sys_pc2epc = _RANDOM[11'h4A8][10];	// rob.scala:310:28
        rob_uop_2_26_flush_on_commit = _RANDOM[11'h4A8][12];	// rob.scala:310:28
        rob_uop_2_26_ldst = _RANDOM[11'h4A8][19:14];	// rob.scala:310:28
        rob_uop_2_26_ldst_val = _RANDOM[11'h4A9][6];	// rob.scala:310:28
        rob_uop_2_26_dst_rtype = _RANDOM[11'h4A9][8:7];	// rob.scala:310:28
        rob_uop_2_26_fp_val = _RANDOM[11'h4A9][14];	// rob.scala:310:28
        rob_uop_2_27_uopc = _RANDOM[11'h4A9][31:25];	// rob.scala:310:28
        rob_uop_2_27_is_rvc = _RANDOM[11'h4AC][0];	// rob.scala:310:28
        rob_uop_2_27_br_mask = {_RANDOM[11'h4AE][31:21], _RANDOM[11'h4AF][4:0]};	// rob.scala:310:28
        rob_uop_2_27_ftq_idx = _RANDOM[11'h4AF][13:9];	// rob.scala:310:28
        rob_uop_2_27_edge_inst = _RANDOM[11'h4AF][14];	// rob.scala:310:28
        rob_uop_2_27_pc_lob = _RANDOM[11'h4AF][20:15];	// rob.scala:310:28
        rob_uop_2_27_pdst = _RANDOM[11'h4B1][15:9];	// rob.scala:310:28
        rob_uop_2_27_stale_pdst = _RANDOM[11'h4B2][20:14];	// rob.scala:310:28
        rob_uop_2_27_is_fencei = _RANDOM[11'h4B5][0];	// rob.scala:310:28
        rob_uop_2_27_uses_ldq = _RANDOM[11'h4B5][2];	// rob.scala:310:28
        rob_uop_2_27_uses_stq = _RANDOM[11'h4B5][3];	// rob.scala:310:28
        rob_uop_2_27_is_sys_pc2epc = _RANDOM[11'h4B5][4];	// rob.scala:310:28
        rob_uop_2_27_flush_on_commit = _RANDOM[11'h4B5][6];	// rob.scala:310:28
        rob_uop_2_27_ldst = _RANDOM[11'h4B5][13:8];	// rob.scala:310:28
        rob_uop_2_27_ldst_val = _RANDOM[11'h4B6][0];	// rob.scala:310:28
        rob_uop_2_27_dst_rtype = _RANDOM[11'h4B6][2:1];	// rob.scala:310:28
        rob_uop_2_27_fp_val = _RANDOM[11'h4B6][8];	// rob.scala:310:28
        rob_uop_2_28_uopc = _RANDOM[11'h4B6][25:19];	// rob.scala:310:28
        rob_uop_2_28_is_rvc = _RANDOM[11'h4B8][26];	// rob.scala:310:28
        rob_uop_2_28_br_mask = _RANDOM[11'h4BB][30:15];	// rob.scala:310:28
        rob_uop_2_28_ftq_idx = _RANDOM[11'h4BC][7:3];	// rob.scala:310:28
        rob_uop_2_28_edge_inst = _RANDOM[11'h4BC][8];	// rob.scala:310:28
        rob_uop_2_28_pc_lob = _RANDOM[11'h4BC][14:9];	// rob.scala:310:28
        rob_uop_2_28_pdst = _RANDOM[11'h4BE][9:3];	// rob.scala:310:28
        rob_uop_2_28_stale_pdst = _RANDOM[11'h4BF][14:8];	// rob.scala:310:28
        rob_uop_2_28_is_fencei = _RANDOM[11'h4C1][26];	// rob.scala:310:28
        rob_uop_2_28_uses_ldq = _RANDOM[11'h4C1][28];	// rob.scala:310:28
        rob_uop_2_28_uses_stq = _RANDOM[11'h4C1][29];	// rob.scala:310:28
        rob_uop_2_28_is_sys_pc2epc = _RANDOM[11'h4C1][30];	// rob.scala:310:28
        rob_uop_2_28_flush_on_commit = _RANDOM[11'h4C2][0];	// rob.scala:310:28
        rob_uop_2_28_ldst = _RANDOM[11'h4C2][7:2];	// rob.scala:310:28
        rob_uop_2_28_ldst_val = _RANDOM[11'h4C2][26];	// rob.scala:310:28
        rob_uop_2_28_dst_rtype = _RANDOM[11'h4C2][28:27];	// rob.scala:310:28
        rob_uop_2_28_fp_val = _RANDOM[11'h4C3][2];	// rob.scala:310:28
        rob_uop_2_29_uopc = _RANDOM[11'h4C3][19:13];	// rob.scala:310:28
        rob_uop_2_29_is_rvc = _RANDOM[11'h4C5][20];	// rob.scala:310:28
        rob_uop_2_29_br_mask = _RANDOM[11'h4C8][24:9];	// rob.scala:310:28
        rob_uop_2_29_ftq_idx = {_RANDOM[11'h4C8][31:29], _RANDOM[11'h4C9][1:0]};	// rob.scala:310:28
        rob_uop_2_29_edge_inst = _RANDOM[11'h4C9][2];	// rob.scala:310:28
        rob_uop_2_29_pc_lob = _RANDOM[11'h4C9][8:3];	// rob.scala:310:28
        rob_uop_2_29_pdst = {_RANDOM[11'h4CA][31:29], _RANDOM[11'h4CB][3:0]};	// rob.scala:310:28
        rob_uop_2_29_stale_pdst = _RANDOM[11'h4CC][8:2];	// rob.scala:310:28
        rob_uop_2_29_is_fencei = _RANDOM[11'h4CE][20];	// rob.scala:310:28
        rob_uop_2_29_uses_ldq = _RANDOM[11'h4CE][22];	// rob.scala:310:28
        rob_uop_2_29_uses_stq = _RANDOM[11'h4CE][23];	// rob.scala:310:28
        rob_uop_2_29_is_sys_pc2epc = _RANDOM[11'h4CE][24];	// rob.scala:310:28
        rob_uop_2_29_flush_on_commit = _RANDOM[11'h4CE][26];	// rob.scala:310:28
        rob_uop_2_29_ldst = {_RANDOM[11'h4CE][31:28], _RANDOM[11'h4CF][1:0]};	// rob.scala:310:28
        rob_uop_2_29_ldst_val = _RANDOM[11'h4CF][20];	// rob.scala:310:28
        rob_uop_2_29_dst_rtype = _RANDOM[11'h4CF][22:21];	// rob.scala:310:28
        rob_uop_2_29_fp_val = _RANDOM[11'h4CF][28];	// rob.scala:310:28
        rob_uop_2_30_uopc = _RANDOM[11'h4D0][13:7];	// rob.scala:310:28
        rob_uop_2_30_is_rvc = _RANDOM[11'h4D2][14];	// rob.scala:310:28
        rob_uop_2_30_br_mask = _RANDOM[11'h4D5][18:3];	// rob.scala:310:28
        rob_uop_2_30_ftq_idx = _RANDOM[11'h4D5][27:23];	// rob.scala:310:28
        rob_uop_2_30_edge_inst = _RANDOM[11'h4D5][28];	// rob.scala:310:28
        rob_uop_2_30_pc_lob = {_RANDOM[11'h4D5][31:29], _RANDOM[11'h4D6][2:0]};	// rob.scala:310:28
        rob_uop_2_30_pdst = _RANDOM[11'h4D7][29:23];	// rob.scala:310:28
        rob_uop_2_30_stale_pdst = {_RANDOM[11'h4D8][31:28], _RANDOM[11'h4D9][2:0]};	// rob.scala:310:28
        rob_uop_2_30_is_fencei = _RANDOM[11'h4DB][14];	// rob.scala:310:28
        rob_uop_2_30_uses_ldq = _RANDOM[11'h4DB][16];	// rob.scala:310:28
        rob_uop_2_30_uses_stq = _RANDOM[11'h4DB][17];	// rob.scala:310:28
        rob_uop_2_30_is_sys_pc2epc = _RANDOM[11'h4DB][18];	// rob.scala:310:28
        rob_uop_2_30_flush_on_commit = _RANDOM[11'h4DB][20];	// rob.scala:310:28
        rob_uop_2_30_ldst = _RANDOM[11'h4DB][27:22];	// rob.scala:310:28
        rob_uop_2_30_ldst_val = _RANDOM[11'h4DC][14];	// rob.scala:310:28
        rob_uop_2_30_dst_rtype = _RANDOM[11'h4DC][16:15];	// rob.scala:310:28
        rob_uop_2_30_fp_val = _RANDOM[11'h4DC][22];	// rob.scala:310:28
        rob_uop_2_31_uopc = _RANDOM[11'h4DD][7:1];	// rob.scala:310:28
        rob_uop_2_31_is_rvc = _RANDOM[11'h4DF][8];	// rob.scala:310:28
        rob_uop_2_31_br_mask = {_RANDOM[11'h4E1][31:29], _RANDOM[11'h4E2][12:0]};	// rob.scala:310:28
        rob_uop_2_31_ftq_idx = _RANDOM[11'h4E2][21:17];	// rob.scala:310:28
        rob_uop_2_31_edge_inst = _RANDOM[11'h4E2][22];	// rob.scala:310:28
        rob_uop_2_31_pc_lob = _RANDOM[11'h4E2][28:23];	// rob.scala:310:28
        rob_uop_2_31_pdst = _RANDOM[11'h4E4][23:17];	// rob.scala:310:28
        rob_uop_2_31_stale_pdst = _RANDOM[11'h4E5][28:22];	// rob.scala:310:28
        rob_uop_2_31_is_fencei = _RANDOM[11'h4E8][8];	// rob.scala:310:28
        rob_uop_2_31_uses_ldq = _RANDOM[11'h4E8][10];	// rob.scala:310:28
        rob_uop_2_31_uses_stq = _RANDOM[11'h4E8][11];	// rob.scala:310:28
        rob_uop_2_31_is_sys_pc2epc = _RANDOM[11'h4E8][12];	// rob.scala:310:28
        rob_uop_2_31_flush_on_commit = _RANDOM[11'h4E8][14];	// rob.scala:310:28
        rob_uop_2_31_ldst = _RANDOM[11'h4E8][21:16];	// rob.scala:310:28
        rob_uop_2_31_ldst_val = _RANDOM[11'h4E9][8];	// rob.scala:310:28
        rob_uop_2_31_dst_rtype = _RANDOM[11'h4E9][10:9];	// rob.scala:310:28
        rob_uop_2_31_fp_val = _RANDOM[11'h4E9][16];	// rob.scala:310:28
        rob_exception_2_0 = _RANDOM[11'h4E9][27];	// rob.scala:310:28, :311:28
        rob_exception_2_1 = _RANDOM[11'h4E9][28];	// rob.scala:310:28, :311:28
        rob_exception_2_2 = _RANDOM[11'h4E9][29];	// rob.scala:310:28, :311:28
        rob_exception_2_3 = _RANDOM[11'h4E9][30];	// rob.scala:310:28, :311:28
        rob_exception_2_4 = _RANDOM[11'h4E9][31];	// rob.scala:310:28, :311:28
        rob_exception_2_5 = _RANDOM[11'h4EA][0];	// rob.scala:311:28
        rob_exception_2_6 = _RANDOM[11'h4EA][1];	// rob.scala:311:28
        rob_exception_2_7 = _RANDOM[11'h4EA][2];	// rob.scala:311:28
        rob_exception_2_8 = _RANDOM[11'h4EA][3];	// rob.scala:311:28
        rob_exception_2_9 = _RANDOM[11'h4EA][4];	// rob.scala:311:28
        rob_exception_2_10 = _RANDOM[11'h4EA][5];	// rob.scala:311:28
        rob_exception_2_11 = _RANDOM[11'h4EA][6];	// rob.scala:311:28
        rob_exception_2_12 = _RANDOM[11'h4EA][7];	// rob.scala:311:28
        rob_exception_2_13 = _RANDOM[11'h4EA][8];	// rob.scala:311:28
        rob_exception_2_14 = _RANDOM[11'h4EA][9];	// rob.scala:311:28
        rob_exception_2_15 = _RANDOM[11'h4EA][10];	// rob.scala:311:28
        rob_exception_2_16 = _RANDOM[11'h4EA][11];	// rob.scala:311:28
        rob_exception_2_17 = _RANDOM[11'h4EA][12];	// rob.scala:311:28
        rob_exception_2_18 = _RANDOM[11'h4EA][13];	// rob.scala:311:28
        rob_exception_2_19 = _RANDOM[11'h4EA][14];	// rob.scala:311:28
        rob_exception_2_20 = _RANDOM[11'h4EA][15];	// rob.scala:311:28
        rob_exception_2_21 = _RANDOM[11'h4EA][16];	// rob.scala:311:28
        rob_exception_2_22 = _RANDOM[11'h4EA][17];	// rob.scala:311:28
        rob_exception_2_23 = _RANDOM[11'h4EA][18];	// rob.scala:311:28
        rob_exception_2_24 = _RANDOM[11'h4EA][19];	// rob.scala:311:28
        rob_exception_2_25 = _RANDOM[11'h4EA][20];	// rob.scala:311:28
        rob_exception_2_26 = _RANDOM[11'h4EA][21];	// rob.scala:311:28
        rob_exception_2_27 = _RANDOM[11'h4EA][22];	// rob.scala:311:28
        rob_exception_2_28 = _RANDOM[11'h4EA][23];	// rob.scala:311:28
        rob_exception_2_29 = _RANDOM[11'h4EA][24];	// rob.scala:311:28
        rob_exception_2_30 = _RANDOM[11'h4EA][25];	// rob.scala:311:28
        rob_exception_2_31 = _RANDOM[11'h4EA][26];	// rob.scala:311:28
        rob_predicated_2_0 = _RANDOM[11'h4EA][27];	// rob.scala:311:28, :312:29
        rob_predicated_2_1 = _RANDOM[11'h4EA][28];	// rob.scala:311:28, :312:29
        rob_predicated_2_2 = _RANDOM[11'h4EA][29];	// rob.scala:311:28, :312:29
        rob_predicated_2_3 = _RANDOM[11'h4EA][30];	// rob.scala:311:28, :312:29
        rob_predicated_2_4 = _RANDOM[11'h4EA][31];	// rob.scala:311:28, :312:29
        rob_predicated_2_5 = _RANDOM[11'h4EB][0];	// rob.scala:312:29
        rob_predicated_2_6 = _RANDOM[11'h4EB][1];	// rob.scala:312:29
        rob_predicated_2_7 = _RANDOM[11'h4EB][2];	// rob.scala:312:29
        rob_predicated_2_8 = _RANDOM[11'h4EB][3];	// rob.scala:312:29
        rob_predicated_2_9 = _RANDOM[11'h4EB][4];	// rob.scala:312:29
        rob_predicated_2_10 = _RANDOM[11'h4EB][5];	// rob.scala:312:29
        rob_predicated_2_11 = _RANDOM[11'h4EB][6];	// rob.scala:312:29
        rob_predicated_2_12 = _RANDOM[11'h4EB][7];	// rob.scala:312:29
        rob_predicated_2_13 = _RANDOM[11'h4EB][8];	// rob.scala:312:29
        rob_predicated_2_14 = _RANDOM[11'h4EB][9];	// rob.scala:312:29
        rob_predicated_2_15 = _RANDOM[11'h4EB][10];	// rob.scala:312:29
        rob_predicated_2_16 = _RANDOM[11'h4EB][11];	// rob.scala:312:29
        rob_predicated_2_17 = _RANDOM[11'h4EB][12];	// rob.scala:312:29
        rob_predicated_2_18 = _RANDOM[11'h4EB][13];	// rob.scala:312:29
        rob_predicated_2_19 = _RANDOM[11'h4EB][14];	// rob.scala:312:29
        rob_predicated_2_20 = _RANDOM[11'h4EB][15];	// rob.scala:312:29
        rob_predicated_2_21 = _RANDOM[11'h4EB][16];	// rob.scala:312:29
        rob_predicated_2_22 = _RANDOM[11'h4EB][17];	// rob.scala:312:29
        rob_predicated_2_23 = _RANDOM[11'h4EB][18];	// rob.scala:312:29
        rob_predicated_2_24 = _RANDOM[11'h4EB][19];	// rob.scala:312:29
        rob_predicated_2_25 = _RANDOM[11'h4EB][20];	// rob.scala:312:29
        rob_predicated_2_26 = _RANDOM[11'h4EB][21];	// rob.scala:312:29
        rob_predicated_2_27 = _RANDOM[11'h4EB][22];	// rob.scala:312:29
        rob_predicated_2_28 = _RANDOM[11'h4EB][23];	// rob.scala:312:29
        rob_predicated_2_29 = _RANDOM[11'h4EB][24];	// rob.scala:312:29
        rob_predicated_2_30 = _RANDOM[11'h4EB][25];	// rob.scala:312:29
        rob_predicated_2_31 = _RANDOM[11'h4EB][26];	// rob.scala:312:29
        block_commit_REG = _RANDOM[11'h4EB][27];	// rob.scala:312:29, :540:94
        block_commit_REG_1 = _RANDOM[11'h4EB][28];	// rob.scala:312:29, :540:131
        block_commit_REG_2 = _RANDOM[11'h4EB][29];	// rob.scala:312:29, :540:123
        r_partial_row = _RANDOM[11'h4EB][30];	// rob.scala:312:29, :677:30
        pnr_maybe_at_tail = _RANDOM[11'h4EB][31];	// rob.scala:312:29, :714:36
        REG = _RANDOM[11'h4EC][0];	// rob.scala:808:30
        REG_1 = _RANDOM[11'h4EC][1];	// rob.scala:808:{22,30}
        REG_2 = _RANDOM[11'h4EC][2];	// rob.scala:808:30, :824:22
        io_com_load_is_at_rob_head_REG = _RANDOM[11'h4EC][3];	// rob.scala:808:30, :865:40
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  rob_fflags_32x5_0 rob_fflags_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_1_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_1_valid & io_fflags_1_bits_uop_rob_idx[1:0] == 2'h0),	// rob.scala:221:26, :272:36, :304:53, :381:32
    .W0_clk  (clock),
    .W0_data (io_fflags_1_bits_flags),
    .W1_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h0),	// rob.scala:221:26, :272:36, :304:53, :381:32
    .W1_clk  (clock),
    .W1_data (io_fflags_0_bits_flags),
    .W2_addr (rob_tail),	// rob.scala:228:29
    .W2_en   (io_enq_valids_0),
    .W2_clk  (clock),
    .W2_data (5'h0),	// rob.scala:224:29
    .R0_data (_rob_fflags_ext_R0_data)
  );
  rob_fflags_32x5_0 rob_fflags_1_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_1_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_1_valid & io_fflags_1_bits_uop_rob_idx[1:0] == 2'h1),	// rob.scala:272:36, :304:53, :381:32, :540:33
    .W0_clk  (clock),
    .W0_data (io_fflags_1_bits_flags),
    .W1_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h1),	// rob.scala:272:36, :304:53, :381:32, :540:33
    .W1_clk  (clock),
    .W1_data (io_fflags_0_bits_flags),
    .W2_addr (rob_tail),	// rob.scala:228:29
    .W2_en   (io_enq_valids_1),
    .W2_clk  (clock),
    .W2_data (5'h0),	// rob.scala:224:29
    .R0_data (_rob_fflags_1_ext_R0_data)
  );
  rob_fflags_32x5_0 rob_fflags_2_ext (	// rob.scala:313:28
    .R0_addr (rob_head),	// rob.scala:224:29
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .W0_addr (io_fflags_1_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W0_en   (io_fflags_1_valid & io_fflags_1_bits_uop_rob_idx[1:0] == 2'h2),	// rob.scala:236:31, :272:36, :304:53, :381:32
    .W0_clk  (clock),
    .W0_data (io_fflags_1_bits_flags),
    .W1_addr (io_fflags_0_bits_uop_rob_idx[6:2]),	// rob.scala:236:31, :268:25
    .W1_en   (io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h2),	// rob.scala:236:31, :272:36, :304:53, :381:32
    .W1_clk  (clock),
    .W1_data (io_fflags_0_bits_flags),
    .W2_addr (rob_tail),	// rob.scala:228:29
    .W2_en   (io_enq_valids_2),
    .W2_clk  (clock),
    .W2_data (5'h0),	// rob.scala:224:29
    .R0_data (_rob_fflags_2_ext_R0_data)
  );
  assign io_rob_tail_idx = rob_tail_idx;	// Cat.scala:30:58
  assign io_rob_head_idx = rob_head_idx;	// Cat.scala:30:58
  assign io_commit_valids_0 = will_commit_0;	// rob.scala:547:70
  assign io_commit_valids_1 = will_commit_1;	// rob.scala:547:70
  assign io_commit_valids_2 = will_commit_2;	// rob.scala:547:70
  assign io_commit_arch_valids_0 = will_commit_0 & ~_GEN_12[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_arch_valids_1 = will_commit_1 & ~_GEN_42[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_arch_valids_2 = will_commit_2 & ~_GEN_72[com_idx];	// rob.scala:236:20, :410:{48,51}, :547:70
  assign io_commit_uops_0_ftq_idx = _GEN_15[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_pdst = _GEN_18[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_stale_pdst = _GEN_19[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_is_fencei = _GEN_20[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_uses_ldq = _GEN_21[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_uses_stq = _GEN_22[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_ldst = _GEN_25[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_ldst_val = _GEN_26[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_0_dst_rtype = _GEN_27[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_ftq_idx = _GEN_45[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_pdst = _GEN_48[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_stale_pdst = _GEN_49[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_is_fencei = _GEN_50[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_uses_ldq = _GEN_51[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_uses_stq = _GEN_52[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_ldst = _GEN_55[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_ldst_val = _GEN_56[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_1_dst_rtype = _GEN_57[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_ftq_idx = _GEN_75[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_pdst = _GEN_78[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_stale_pdst = _GEN_79[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_is_fencei = _GEN_80[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_uses_ldq = _GEN_81[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_uses_stq = _GEN_82[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_ldst = _GEN_85[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_ldst_val = _GEN_86[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_uops_2_dst_rtype = _GEN_87[com_idx];	// rob.scala:236:20, :411:25
  assign io_commit_fflags_valid = fflags_val_0 | fflags_val_1 | fflags_val_2;	// rob.scala:602:32, :617:48
  assign io_commit_fflags_bits =
    (fflags_val_0 ? _rob_fflags_ext_R0_data : 5'h0)
    | (fflags_val_1 ? _rob_fflags_1_ext_R0_data : 5'h0)
    | (fflags_val_2 ? _rob_fflags_2_ext_R0_data : 5'h0);	// rob.scala:224:29, :313:28, :602:32, :605:21, :618:44
  assign io_commit_rbk_valids_0 = _io_commit_rbk_valids_0_output;	// rob.scala:427:40
  assign io_commit_rbk_valids_1 = _io_commit_rbk_valids_1_output;	// rob.scala:427:40
  assign io_commit_rbk_valids_2 = _io_commit_rbk_valids_2_output;	// rob.scala:427:40
  assign io_commit_rollback = _io_commit_rollback_T_2;	// rob.scala:236:31
  assign io_com_load_is_at_rob_head = io_com_load_is_at_rob_head_REG;	// rob.scala:865:40
  assign io_com_xcpt_valid = exception_thrown & _io_flush_bits_flush_typ_T;	// rob.scala:545:85, :556:50, :557:41
  assign io_com_xcpt_bits_ftq_idx = com_xcpt_uop_ftq_idx;	// Mux.scala:47:69
  assign io_com_xcpt_bits_edge_inst = com_xcpt_uop_edge_inst;	// Mux.scala:47:69
  assign io_com_xcpt_bits_pc_lob = com_xcpt_uop_pc_lob;	// Mux.scala:47:69
  assign io_com_xcpt_bits_cause = r_xcpt_uop_exc_cause;	// rob.scala:259:29
  assign io_com_xcpt_bits_badvaddr = {{24{r_xcpt_badvaddr[39]}}, r_xcpt_badvaddr};	// Bitwise.scala:72:12, Cat.scala:30:58, rob.scala:260:29, util.scala:261:46
  assign io_flush_valid = _io_flush_valid_output;	// rob.scala:573:36
  assign io_flush_bits_ftq_idx =
    exception_thrown
      ? com_xcpt_uop_ftq_idx
      : (flush_commit_mask_0 ? _GEN_15[com_idx] : 5'h0)
        | (flush_commit_mask_1 ? _GEN_45[com_idx] : 5'h0)
        | (flush_commit_mask_2 ? _GEN_75[com_idx] : 5'h0);	// Mux.scala:27:72, :47:69, rob.scala:224:29, :236:20, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_edge_inst =
    exception_thrown
      ? com_xcpt_uop_edge_inst
      : flush_commit_mask_0 & _GEN_16[com_idx] | flush_commit_mask_1 & _GEN_46[com_idx]
        | flush_commit_mask_2 & _GEN_76[com_idx];	// Mux.scala:27:72, :47:69, rob.scala:236:20, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_is_rvc =
    exception_thrown
      ? (rob_head_vals_0
           ? _GEN_14[com_idx]
           : rob_head_vals_1 ? _GEN_44[com_idx] : _GEN_74[com_idx])
      : flush_commit_mask_0 & _GEN_14[com_idx] | flush_commit_mask_1 & _GEN_44[com_idx]
        | flush_commit_mask_2 & _GEN_74[com_idx];	// Mux.scala:27:72, :47:69, rob.scala:236:20, :398:49, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_pc_lob =
    exception_thrown
      ? com_xcpt_uop_pc_lob
      : (flush_commit_mask_0 ? _GEN_17[com_idx] : 6'h0)
        | (flush_commit_mask_1 ? _GEN_47[com_idx] : 6'h0)
        | (flush_commit_mask_2 ? _GEN_77[com_idx] : 6'h0);	// Mux.scala:27:72, :47:69, rob.scala:236:20, :287:15, :411:25, :545:85, :571:75, :578:22
  assign io_flush_bits_flush_typ =
    _io_flush_valid_output
      ? (flush_commit
         & (exception_thrown
              ? (rob_head_vals_0
                   ? _GEN_13[com_idx]
                   : rob_head_vals_1 ? _GEN_43[com_idx] : _GEN_73[com_idx])
              : (flush_commit_mask_0 ? _GEN_13[com_idx] : 7'h0)
                | (flush_commit_mask_1 ? _GEN_43[com_idx] : 7'h0)
                | (flush_commit_mask_2 ? _GEN_73[com_idx] : 7'h0)) == 7'h6A
           ? 3'h3
           : exception_thrown & _io_flush_bits_flush_typ_T
               ? 3'h1
               : exception_thrown | (rob_head_vals_0 | rob_head_vals_1 | rob_head_vals_2)
                 & (rob_head_vals_0
                      ? _GEN_23[com_idx]
                      : rob_head_vals_1 ? _GEN_53[com_idx] : _GEN_83[com_idx])
                   ? 3'h2
                   : 3'h4)
      : 3'h0;	// Mux.scala:27:72, :47:69, rob.scala:172:10, :173:10, :174:10, :175:10, :236:20, :287:15, :398:49, :411:25, :457:33, :545:85, :556:50, :562:{27,31}, :564:39, :571:75, :572:48, :573:36, :578:22, :587:66, :588:{62,80}
  assign io_empty = empty;	// rob.scala:788:41
  assign io_ready = _io_ready_T & ~full & ~r_xcpt_val;	// rob.scala:258:33, :425:47, :658:33, :716:33, :787:39, :794:56
  assign io_flush_frontend = r_xcpt_val;	// rob.scala:258:33
endmodule

